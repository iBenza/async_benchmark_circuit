
module Balsa_gcd8 ( activate_0r, activate_0a, x_0r, x_0a, x_0d, y_0r, y_0a, y_0d, z_0r, z_0a, z_0d, initialise );
  input [7:0] x_0d;
  input [7:0] y_0d;
  output [7:0] z_0d;
  input activate_0r, x_0a, y_0a, z_0a, initialise;
  output activate_0a, x_0r, y_0r, z_0r;

  wire activate_0r;
  wire activate_0a;
  wire x_0r;
  wire x_0a;
  wire [7:0] x_0d;
  wire y_0r;
  wire y_0a;
  wire [7:0] y_0d;
  wire z_0r;
  wire z_0a;
  wire [7:0] z_0d;
  wire initialise;
  wire c45_r;
  wire c45_a;
  wire [7:0] c45_d;
  wire c44_r;
  wire c44_a;
  wire [7:0] c44_d;
  wire c43_r;
  wire c42_r;
  wire c42_a;
  wire c40_a;
  wire c38_a;
  wire c37_r;
  wire c37_a;
  wire c36_r;
  wire c36_a;
  wire c36_d;
  wire [7:0] c34_d;
  wire c33_r;
  wire c33_d;
  wire c32_r;
  wire c32_d;
  wire c31_a;
  wire c30_a;
  wire c28_r;
  wire c27_r;
  wire [7:0] c24_d;
  wire c23_a;
  wire c22_r;
  wire c21_r;
  wire c20_r;
  wire c19_a;
  wire c18_a;
  wire [7:0] c18_d;
  wire [7:0] c15_d;
  wire c14_a;
  wire c13_r;
  wire c12_r;
  wire c11_r;
  wire c10_a;
  wire c9_a;
  wire [7:0] c9_d;
  wire I0_nbWriteReq_0n;
  wire I0_bWriteReq_0n;
  wire I0_nWriteReq_0n;
  wire I2_nbWriteReq_0n;
  wire I2_bWriteReq_0n;
  wire I2_nWriteReq_0n;
  wire I1_nselect_0n;
  wire I1_select_0n;
  wire I3_nselect_0n;
  wire I3_select_0n;
  wire I4_nReq_0n;
  wire I5_sreq_0n_1_;
  wire I5_I3_s;
  wire [1:0] I6_acks_0n;
  wire I6_I1_s_0n;
  wire I6_I2_s_0n;
  wire I9_nReq_0n;
  wire I9_guardAck_0n;
  wire I9_guardReq_0n;
  wire [7:0] I10_eq_0n;
  wire [1:0] I10_internal_0n;
  wire I9_I0_ns_0n;
  wire I11_I5_ns_0n;
  wire I15_nbWriteReq_0n;
  wire I15_bWriteReq_0n;
  wire I15_nWriteReq_0n;
  wire I16_vcc;
  wire I16_nxv_0n;
  wire I16_z_0n;
  wire I16_v_0n;
  wire [7:0] I16_n_0n;
  wire I16_addOut_0n_0_;
  wire I16_addOut_0n_1_;
  wire I16_addOut_0n_2_;
  wire I16_addOut_0n_3_;
  wire I16_addOut_0n_4_;
  wire I16_addOut_0n_5_;
  wire I16_addOut_0n_6_;
  wire I16_addOut_0n_7_;
  wire I16_c_0n_1_;
  wire I16_c_0n_2_;
  wire I16_c_0n_3_;
  wire I16_c_0n_4_;
  wire I16_c_0n_5_;
  wire I16_c_0n_6_;
  wire I16_c_0n_7_;
  wire I16_c_0n_8_;
  wire I16_nCv_0n_1_;
  wire I16_nCv_0n_2_;
  wire I16_nCv_0n_3_;
  wire I16_nCv_0n_4_;
  wire I16_nCv_0n_5_;
  wire I16_nCv_0n_6_;
  wire I16_nCv_0n_7_;
  wire I16_nCv_0n_8_;
  wire I16_nStart_0n;
  wire I16_start_0n;
  wire [3:0] I16_internal_0n;
  wire I5_I4_s_0n;
  wire I9_I1_s_0n;
  wire I12_I3_s_0n;
  wire I17_I3_s_0n;
  wire I22_I3_s_0n;
  wire I20_nbWriteReq_0n;
  wire I20_bWriteReq_0n;
  wire I20_nWriteReq_0n;
  wire I25_nbWriteReq_0n;
  wire I25_bWriteReq_0n;
  wire I25_nWriteReq_0n;
  wire I21_vcc;
  wire [7:0] I21_n_0n;
  wire [8:1] I21_c_0n;
  wire I21_nCv_0n_1_;
  wire I21_nCv_0n_2_;
  wire I21_nCv_0n_3_;
  wire I21_nCv_0n_4_;
  wire I21_nCv_0n_5_;
  wire I21_nCv_0n_6_;
  wire I21_nCv_0n_7_;
  wire I21_nCv_0n_8_;
  wire I21_nStart_0n;
  wire I21_start_0n;
  wire [1:0] I21_internal_0n;
  wire I26_vcc;
  wire [7:0] I26_n_0n;
  wire [8:1] I26_c_0n;
  wire I26_nCv_0n_1_;
  wire I26_nCv_0n_2_;
  wire I26_nCv_0n_3_;
  wire I26_nCv_0n_4_;
  wire I26_nCv_0n_5_;
  wire I26_nCv_0n_6_;
  wire I26_nCv_0n_7_;
  wire I26_nCv_0n_8_;
  wire I26_nStart_0n;
  wire I26_start_0n;
  wire [1:0] I26_internal_0n;
  wire I16_I9_cv;
  wire I16_I9_ha;
  wire I16_I9_start;
  wire I16_I10_cv;
  wire I16_I10_ha;
  wire I16_I10_start;
  wire I16_I11_cv;
  wire I16_I11_ha;
  wire I16_I11_start;
  wire I16_I12_cv;
  wire I16_I12_ha;
  wire I16_I12_start;
  wire I16_I13_cv;
  wire I16_I13_ha;
  wire I16_I13_start;
  wire I16_I14_cv;
  wire I16_I14_ha;
  wire I16_I14_start;
  wire I16_I15_cv;
  wire I16_I15_ha;
  wire I16_I15_start;
  wire I16_I16_cv;
  wire I16_I16_ha;
  wire I16_I16_start;
  wire I21_I11_cv;
  wire I21_I11_ha;
  wire I21_I11_start;
  wire I21_I12_cv;
  wire I21_I12_ha;
  wire I21_I12_start;
  wire I21_I13_cv;
  wire I21_I13_ha;
  wire I21_I13_start;
  wire I21_I14_cv;
  wire I21_I14_ha;
  wire I21_I14_start;
  wire I21_I15_cv;
  wire I21_I15_ha;
  wire I21_I15_start;
  wire I21_I16_cv;
  wire I21_I16_ha;
  wire I21_I16_start;
  wire I21_I17_cv;
  wire I21_I17_ha;
  wire I21_I17_start;
  wire I21_I18_cv;
  wire I21_I18_ha;
  wire I21_I18_start;
  wire I26_I11_cv;
  wire I26_I11_ha;
  wire I26_I11_start;
  wire I26_I12_cv;
  wire I26_I12_ha;
  wire I26_I12_start;
  wire I26_I13_cv;
  wire I26_I13_ha;
  wire I26_I13_start;
  wire I26_I14_cv;
  wire I26_I14_ha;
  wire I26_I14_start;
  wire I26_I15_cv;
  wire I26_I15_ha;
  wire I26_I15_start;
  wire I26_I16_cv;
  wire I26_I16_ha;
  wire I26_I16_start;
  wire I26_I17_cv;
  wire I26_I17_ha;
  wire I26_I17_start;
  wire I26_I18_cv;
  wire I26_I18_ha;
  wire I26_I18_start;
  wire I16_I9_I2_nsel_0n;
  wire I16_I10_I2_nsel_0n;
  wire I16_I11_I2_nsel_0n;
  wire I16_I12_I2_nsel_0n;
  wire I16_I13_I2_nsel_0n;
  wire I16_I14_I2_nsel_0n;
  wire I16_I15_I2_nsel_0n;
  wire I16_I16_I2_nsel_0n;
  wire I21_I11_I2_nsel_0n;
  wire I21_I12_I2_nsel_0n;
  wire I21_I13_I2_nsel_0n;
  wire I21_I14_I2_nsel_0n;
  wire I21_I15_I2_nsel_0n;
  wire I21_I16_I2_nsel_0n;
  wire I21_I17_I2_nsel_0n;
  wire I21_I18_I2_nsel_0n;
  wire I26_I11_I2_nsel_0n;
  wire I26_I12_I2_nsel_0n;
  wire I26_I13_I2_nsel_0n;
  wire I26_I14_I2_nsel_0n;
  wire I26_I15_I2_nsel_0n;
  wire I26_I16_I2_nsel_0n;
  wire I26_I17_I2_nsel_0n;
  wire I26_I18_I2_nsel_0n;
  wire [1:0] I16_I9_I2_I0_int_0n;
  wire [1:0] I16_I10_I2_I0_int_0n;
  wire [1:0] I16_I11_I2_I0_int_0n;
  wire [1:0] I16_I12_I2_I0_int_0n;
  wire [1:0] I16_I13_I2_I0_int_0n;
  wire [1:0] I16_I14_I2_I0_int_0n;
  wire [1:0] I16_I15_I2_I0_int_0n;
  wire [1:0] I16_I16_I2_I0_int_0n;
  wire [1:0] I21_I11_I2_I0_int_0n;
  wire [1:0] I21_I12_I2_I0_int_0n;
  wire [1:0] I21_I13_I2_I0_int_0n;
  wire [1:0] I21_I14_I2_I0_int_0n;
  wire [1:0] I21_I15_I2_I0_int_0n;
  wire [1:0] I21_I16_I2_I0_int_0n;
  wire [1:0] I21_I17_I2_I0_int_0n;
  wire [1:0] I21_I18_I2_I0_int_0n;
  wire [1:0] I26_I11_I2_I0_int_0n;
  wire [1:0] I26_I12_I2_I0_int_0n;
  wire [1:0] I26_I13_I2_I0_int_0n;
  wire [1:0] I26_I14_I2_I0_int_0n;
  wire [1:0] I26_I15_I2_I0_int_0n;
  wire [1:0] I26_I16_I2_I0_int_0n;
  wire [1:0] I26_I17_I2_I0_int_0n;
  wire [1:0] I26_I18_I2_I0_int_0n;
  wire I1_I0_nsel_0n;
  wire I1_I1_nsel_0n;
  wire I1_I2_nsel_0n;
  wire I1_I3_nsel_0n;
  wire I1_I4_nsel_0n;
  wire I1_I5_nsel_0n;
  wire I1_I6_nsel_0n;
  wire I1_I7_nsel_0n;
  wire I1_I8_nsel_0n;
  wire I3_I0_nsel_0n;
  wire I3_I1_nsel_0n;
  wire I3_I2_nsel_0n;
  wire I3_I3_nsel_0n;
  wire I3_I4_nsel_0n;
  wire I3_I5_nsel_0n;
  wire I3_I6_nsel_0n;
  wire I3_I7_nsel_0n;
  wire I3_I8_nsel_0n;
  wire I16_I9_I3_nsel_0n;
  wire I16_I10_I3_nsel_0n;
  wire I16_I11_I3_nsel_0n;
  wire I16_I12_I3_nsel_0n;
  wire I16_I13_I3_nsel_0n;
  wire I16_I14_I3_nsel_0n;
  wire I16_I15_I3_nsel_0n;
  wire I16_I16_I3_nsel_0n;
  wire I21_I11_I3_nsel_0n;
  wire I21_I12_I3_nsel_0n;
  wire I21_I13_I3_nsel_0n;
  wire I21_I14_I3_nsel_0n;
  wire I21_I15_I3_nsel_0n;
  wire I21_I16_I3_nsel_0n;
  wire I21_I17_I3_nsel_0n;
  wire I21_I18_I3_nsel_0n;
  wire I26_I11_I3_nsel_0n;
  wire I26_I12_I3_nsel_0n;
  wire I26_I13_I3_nsel_0n;
  wire I26_I14_I3_nsel_0n;
  wire I26_I15_I3_nsel_0n;
  wire I26_I16_I3_nsel_0n;
  wire I26_I17_I3_nsel_0n;
  wire I26_I18_I3_nsel_0n;
  wire [1:0] I1_I0_I0_int_0n;
  wire [1:0] I1_I1_I0_int_0n;
  wire [1:0] I1_I2_I0_int_0n;
  wire [1:0] I1_I3_I0_int_0n;
  wire [1:0] I1_I4_I0_int_0n;
  wire [1:0] I1_I5_I0_int_0n;
  wire [1:0] I1_I6_I0_int_0n;
  wire [1:0] I1_I7_I0_int_0n;
  wire [1:0] I1_I8_I0_int_0n;
  wire [1:0] I3_I0_I0_int_0n;
  wire [1:0] I3_I1_I0_int_0n;
  wire [1:0] I3_I2_I0_int_0n;
  wire [1:0] I3_I3_I0_int_0n;
  wire [1:0] I3_I4_I0_int_0n;
  wire [1:0] I3_I5_I0_int_0n;
  wire [1:0] I3_I6_I0_int_0n;
  wire [1:0] I3_I7_I0_int_0n;
  wire [1:0] I3_I8_I0_int_0n;
  wire [1:0] I16_I9_I3_I0_int_0n;
  wire [1:0] I16_I10_I3_I0_int_0n;
  wire [1:0] I16_I11_I3_I0_int_0n;
  wire [1:0] I16_I12_I3_I0_int_0n;
  wire [1:0] I16_I13_I3_I0_int_0n;
  wire [1:0] I16_I14_I3_I0_int_0n;
  wire [1:0] I16_I15_I3_I0_int_0n;
  wire [1:0] I16_I16_I3_I0_int_0n;
  wire [1:0] I21_I11_I3_I0_int_0n;
  wire [1:0] I21_I12_I3_I0_int_0n;
  wire [1:0] I21_I13_I3_I0_int_0n;
  wire [1:0] I21_I14_I3_I0_int_0n;
  wire [1:0] I21_I15_I3_I0_int_0n;
  wire [1:0] I21_I16_I3_I0_int_0n;
  wire [1:0] I21_I17_I3_I0_int_0n;
  wire [1:0] I21_I18_I3_I0_int_0n;
  wire [1:0] I26_I11_I3_I0_int_0n;
  wire [1:0] I26_I12_I3_I0_int_0n;
  wire [1:0] I26_I13_I3_I0_int_0n;
  wire [1:0] I26_I14_I3_I0_int_0n;
  wire [1:0] I26_I15_I3_I0_int_0n;
  wire [1:0] I26_I16_I3_I0_int_0n;
  wire [1:0] I26_I17_I3_I0_int_0n;
  wire [1:0] I26_I18_I3_I0_int_0n;

  IV I0_I56 ( I0_nWriteReq_0n, c45_r );
  IV I0_I55 ( I0_bWriteReq_0n, I0_nWriteReq_0n );
  IV I0_I54 ( I0_nbWriteReq_0n, I0_bWriteReq_0n );
  IV I0_I53 ( c45_a, I0_nbWriteReq_0n );
  LD1 I0_I52 ( c45_d[7], I0_bWriteReq_0n, z_0d[7] );
  LD1 I0_I51 ( c45_d[6], I0_bWriteReq_0n, z_0d[6] );
  LD1 I0_I50 ( c45_d[5], I0_bWriteReq_0n, z_0d[5] );
  LD1 I0_I49 ( c45_d[4], I0_bWriteReq_0n, z_0d[4] );
  LD1 I0_I48 ( c45_d[3], I0_bWriteReq_0n, z_0d[3] );
  LD1 I0_I47 ( c45_d[2], I0_bWriteReq_0n, z_0d[2] );
  LD1 I0_I46 ( c45_d[1], I0_bWriteReq_0n, z_0d[1] );
  LD1 I0_I45 ( c45_d[0], I0_bWriteReq_0n, z_0d[0] );
  IV I2_I47 ( I2_nWriteReq_0n, c44_r );
  IV I2_I46 ( I2_bWriteReq_0n, I2_nWriteReq_0n );
  IV I2_I45 ( I2_nbWriteReq_0n, I2_bWriteReq_0n );
  IV I2_I44 ( c44_a, I2_nbWriteReq_0n );
  LD1 I2_I43 ( c44_d[7], I2_bWriteReq_0n, c34_d[7] );
  LD1 I2_I42 ( c44_d[6], I2_bWriteReq_0n, c34_d[6] );
  LD1 I2_I41 ( c44_d[5], I2_bWriteReq_0n, c34_d[5] );
  LD1 I2_I40 ( c44_d[4], I2_bWriteReq_0n, c34_d[4] );
  LD1 I2_I39 ( c44_d[3], I2_bWriteReq_0n, c34_d[3] );
  LD1 I2_I38 ( c44_d[2], I2_bWriteReq_0n, c34_d[2] );
  LD1 I2_I37 ( c44_d[1], I2_bWriteReq_0n, c34_d[1] );
  LD1 I2_I36 ( c44_d[0], I2_bWriteReq_0n, c34_d[0] );
  SRFF I1_I11 ( x_0a, c22_r, I1_select_0n, I1_nselect_0n );
  AN2 I1_I10 ( c40_a, I1_select_0n, c45_a );
  AN2 I1_I9 ( c19_a, I1_nselect_0n, c45_a );
  SRFF I3_I11 ( y_0a, c13_r, I3_select_0n, I3_nselect_0n );
  AN2 I3_I10 ( c38_a, I3_select_0n, c44_a );
  AN2 I3_I9 ( c10_a, I3_nselect_0n, c44_a );
  NR2 I4_I1 ( c43_r, I4_nReq_0n, z_0a );
  IV I4_I0 ( I4_nReq_0n, activate_0r );
  GND I4_gnd_cell_instance ( activate_0a );
  C2R I5_I3_I2 ( z_0r, c37_a, I5_sreq_0n_1_, initialise );
  IV I5_I3_I1 ( I5_I3_s, z_0r );
  AN2 I5_I3_I0 ( c37_r, I5_sreq_0n_1_, I5_I3_s );
  C2 I6_I0 ( c42_a, I6_acks_0n[0], I6_acks_0n[1] );
  AN2 I6_I1_I2 ( x_0r, c42_r, I6_I1_s_0n );
  IV I6_I1_I1 ( I6_I1_s_0n, I6_acks_0n[0] );
  ACU0D1 I6_I1_I0 ( I6_acks_0n[0], c40_a, c42_r );
  AN2 I6_I2_I2 ( y_0r, c42_r, I6_I2_s_0n );
  IV I6_I2_I1 ( I6_I2_s_0n, I6_acks_0n[1] );
  ACU0D1 I6_I2_I0 ( I6_acks_0n[1], c38_a, c42_r );
  NR2 I9_I3 ( I9_guardReq_0n, I9_nReq_0n, c31_a );
  IV I9_I2 ( I9_nReq_0n, c37_r );
  C2 I10_I29 ( c36_a, c36_r, c36_r );
  EO I10_I10 ( I10_eq_0n[7], z_0d[7], c34_d[7] );
  EO I10_I9 ( I10_eq_0n[6], z_0d[6], c34_d[6] );
  EO I10_I8 ( I10_eq_0n[5], z_0d[5], c34_d[5] );
  EO I10_I7 ( I10_eq_0n[4], z_0d[4], c34_d[4] );
  EO I10_I6 ( I10_eq_0n[3], z_0d[3], c34_d[3] );
  EO I10_I5 ( I10_eq_0n[2], z_0d[2], c34_d[2] );
  EO I10_I4 ( I10_eq_0n[1], z_0d[1], c34_d[1] );
  EO I10_I3 ( I10_eq_0n[0], z_0d[0], c34_d[0] );
  ND2 I10_I2 ( c36_d, I10_internal_0n[0], I10_internal_0n[1] );
  NR4 I10_I1 ( I10_internal_0n[1], I10_eq_0n[4], I10_eq_0n[5], I10_eq_0n[6], I10_eq_0n[7] );
  NR4 I10_I0 ( I10_internal_0n[0], I10_eq_0n[0], I10_eq_0n[1], I10_eq_0n[2], I10_eq_0n[3] );
  OR2 I11_I0 ( c31_a, c10_a, c19_a );
  IV I9_I0_I2 ( I9_I0_ns_0n, c36_d );
  AN2 I9_I0_I1 ( c37_a, c36_a, I9_I0_ns_0n );
  AN2 I9_I0_I0 ( I9_guardAck_0n, c36_a, c36_d );
  IV I11_I5_I2 ( I11_I5_ns_0n, c33_d );
  AN2 I11_I5_I1 ( c11_r, c33_r, I11_I5_ns_0n );
  AN2 I11_I5_I0 ( c20_r, c33_r, c33_d );
  IV I15_I6 ( I15_nWriteReq_0n, c32_r );
  IV I15_I5 ( I15_bWriteReq_0n, I15_nWriteReq_0n );
  IV I15_I4 ( I15_nbWriteReq_0n, I15_bWriteReq_0n );
  IV I15_I3 ( c30_a, I15_nbWriteReq_0n );
  LD1 I15_I2 ( c32_d, I15_bWriteReq_0n, c33_d );
  C2 I16_I37 ( I16_start_0n, c27_r, c27_r );
  IV I16_I27 ( I16_n_0n[7], c34_d[7] );
  IV I16_I26 ( I16_n_0n[6], c34_d[6] );
  IV I16_I25 ( I16_n_0n[5], c34_d[5] );
  IV I16_I24 ( I16_n_0n[4], c34_d[4] );
  IV I16_I23 ( I16_n_0n[3], c34_d[3] );
  IV I16_I22 ( I16_n_0n[2], c34_d[2] );
  IV I16_I21 ( I16_n_0n[1], c34_d[1] );
  IV I16_I20 ( I16_n_0n[0], c34_d[0] );
  IV I16_I19 ( I16_nStart_0n, I16_start_0n );
  EO I16_I8 ( I16_v_0n, I16_c_0n_7_, I16_c_0n_8_ );
  AN2 I16_I7 ( c32_r, I16_internal_0n[2], I16_internal_0n[3] );
  NR4 I16_I6 ( I16_internal_0n[3], I16_nCv_0n_5_, I16_nCv_0n_6_, I16_nCv_0n_7_, I16_nCv_0n_8_ );
  NR4 I16_I5 ( I16_internal_0n[2], I16_nCv_0n_1_, I16_nCv_0n_2_, I16_nCv_0n_3_, I16_nCv_0n_4_ );
  AN2 I16_I4 ( I16_z_0n, I16_internal_0n[0], I16_internal_0n[1] );
  NR4 I16_I3 ( I16_internal_0n[1], I16_addOut_0n_4_, I16_addOut_0n_5_, I16_addOut_0n_6_, I16_addOut_0n_7_ );
  NR4 I16_I2 ( I16_internal_0n[0], I16_addOut_0n_0_, I16_addOut_0n_1_, I16_addOut_0n_2_, I16_addOut_0n_3_ );
  EO I16_I1 ( I16_nxv_0n, I16_v_0n, I16_addOut_0n_7_ );
  NR2 I16_I0 ( c32_d, I16_z_0n, I16_nxv_0n );
  VCC I16_vcc_cell_instance ( I16_vcc );
  AN2 I5_I4_I2 ( c42_r, c43_r, I5_I4_s_0n );
  NR2 I5_I4_I1 ( I5_sreq_0n_1_, c42_a, I5_I4_s_0n );
  NC2P I5_I4_I0 ( I5_I4_s_0n, c43_r, c42_a );
  AN2 I9_I1_I2 ( c36_r, I9_guardReq_0n, I9_I1_s_0n );
  NR2 I9_I1_I1 ( c28_r, I9_guardAck_0n, I9_I1_s_0n );
  NC2P I9_I1_I0 ( I9_I1_s_0n, I9_guardReq_0n, I9_guardAck_0n );
  AN2 I12_I3_I2 ( c27_r, c28_r, I12_I3_s_0n );
  NR2 I12_I3_I1 ( c33_r, c30_a, I12_I3_s_0n );
  NC2P I12_I3_I0 ( I12_I3_s_0n, c28_r, c30_a );
  AN2 I17_I3_I2 ( c21_r, c20_r, I17_I3_s_0n );
  NR2 I17_I3_I1 ( c22_r, c23_a, I17_I3_s_0n );
  NC2P I17_I3_I0 ( I17_I3_s_0n, c20_r, c23_a );
  AN2 I22_I3_I2 ( c12_r, c11_r, I22_I3_s_0n );
  NR2 I22_I3_I1 ( c13_r, c14_a, I22_I3_s_0n );
  NC2P I22_I3_I0 ( I22_I3_s_0n, c11_r, c14_a );
  IV I20_I20 ( I20_nWriteReq_0n, c18_a );
  IV I20_I19 ( I20_bWriteReq_0n, I20_nWriteReq_0n );
  IV I20_I18 ( I20_nbWriteReq_0n, I20_bWriteReq_0n );
  IV I20_I17 ( c23_a, I20_nbWriteReq_0n );
  LD1 I20_I16 ( c18_d[7], I20_bWriteReq_0n, c24_d[7] );
  LD1 I20_I15 ( c18_d[6], I20_bWriteReq_0n, c24_d[6] );
  LD1 I20_I14 ( c18_d[5], I20_bWriteReq_0n, c24_d[5] );
  LD1 I20_I13 ( c18_d[4], I20_bWriteReq_0n, c24_d[4] );
  LD1 I20_I12 ( c18_d[3], I20_bWriteReq_0n, c24_d[3] );
  LD1 I20_I11 ( c18_d[2], I20_bWriteReq_0n, c24_d[2] );
  LD1 I20_I10 ( c18_d[1], I20_bWriteReq_0n, c24_d[1] );
  LD1 I20_I9 ( c18_d[0], I20_bWriteReq_0n, c24_d[0] );
  IV I25_I20 ( I25_nWriteReq_0n, c9_a );
  IV I25_I19 ( I25_bWriteReq_0n, I25_nWriteReq_0n );
  IV I25_I18 ( I25_nbWriteReq_0n, I25_bWriteReq_0n );
  IV I25_I17 ( c14_a, I25_nbWriteReq_0n );
  LD1 I25_I16 ( c9_d[7], I25_bWriteReq_0n, c15_d[7] );
  LD1 I25_I15 ( c9_d[6], I25_bWriteReq_0n, c15_d[6] );
  LD1 I25_I14 ( c9_d[5], I25_bWriteReq_0n, c15_d[5] );
  LD1 I25_I13 ( c9_d[4], I25_bWriteReq_0n, c15_d[4] );
  LD1 I25_I12 ( c9_d[3], I25_bWriteReq_0n, c15_d[3] );
  LD1 I25_I11 ( c9_d[2], I25_bWriteReq_0n, c15_d[2] );
  LD1 I25_I10 ( c9_d[1], I25_bWriteReq_0n, c15_d[1] );
  LD1 I25_I9 ( c9_d[0], I25_bWriteReq_0n, c15_d[0] );
  C2 I21_I39 ( I21_start_0n, c21_r, c21_r );
  IV I21_I29 ( I21_n_0n[7], c34_d[7] );
  IV I21_I28 ( I21_n_0n[6], c34_d[6] );
  IV I21_I27 ( I21_n_0n[5], c34_d[5] );
  IV I21_I26 ( I21_n_0n[4], c34_d[4] );
  IV I21_I25 ( I21_n_0n[3], c34_d[3] );
  IV I21_I24 ( I21_n_0n[2], c34_d[2] );
  IV I21_I23 ( I21_n_0n[1], c34_d[1] );
  IV I21_I22 ( I21_n_0n[0], c34_d[0] );
  IV I21_I21 ( I21_nStart_0n, I21_start_0n );
  AN2 I21_I2 ( c18_a, I21_internal_0n[0], I21_internal_0n[1] );
  NR4 I21_I1 ( I21_internal_0n[1], I21_nCv_0n_5_, I21_nCv_0n_6_, I21_nCv_0n_7_, I21_nCv_0n_8_ );
  NR4 I21_I0 ( I21_internal_0n[0], I21_nCv_0n_1_, I21_nCv_0n_2_, I21_nCv_0n_3_, I21_nCv_0n_4_ );
  VCC I21_vcc_cell_instance ( I21_vcc );
  C2 I26_I39 ( I26_start_0n, c12_r, c12_r );
  IV I26_I29 ( I26_n_0n[7], z_0d[7] );
  IV I26_I28 ( I26_n_0n[6], z_0d[6] );
  IV I26_I27 ( I26_n_0n[5], z_0d[5] );
  IV I26_I26 ( I26_n_0n[4], z_0d[4] );
  IV I26_I25 ( I26_n_0n[3], z_0d[3] );
  IV I26_I24 ( I26_n_0n[2], z_0d[2] );
  IV I26_I23 ( I26_n_0n[1], z_0d[1] );
  IV I26_I22 ( I26_n_0n[0], z_0d[0] );
  IV I26_I21 ( I26_nStart_0n, I26_start_0n );
  AN2 I26_I2 ( c9_a, I26_internal_0n[0], I26_internal_0n[1] );
  NR4 I26_I1 ( I26_internal_0n[1], I26_nCv_0n_5_, I26_nCv_0n_6_, I26_nCv_0n_7_, I26_nCv_0n_8_ );
  NR4 I26_I0 ( I26_internal_0n[0], I26_nCv_0n_1_, I26_nCv_0n_2_, I26_nCv_0n_3_, I26_nCv_0n_4_ );
  VCC I26_vcc_cell_instance ( I26_vcc );
  EO I16_I9_I5 ( I16_addOut_0n_0_, I16_I9_ha, I16_vcc );
  EO I16_I9_I4 ( I16_I9_ha, I16_n_0n[0], z_0d[0] );
  NR2 I16_I9_I1 ( I16_I9_cv, I16_nStart_0n, I16_nStart_0n );
  IV I16_I9_I0 ( I16_I9_start, I16_nStart_0n );
  EO I16_I10_I5 ( I16_addOut_0n_1_, I16_I10_ha, I16_c_0n_1_ );
  EO I16_I10_I4 ( I16_I10_ha, I16_n_0n[1], z_0d[1] );
  NR2 I16_I10_I1 ( I16_I10_cv, I16_nStart_0n, I16_nCv_0n_1_ );
  IV I16_I10_I0 ( I16_I10_start, I16_nStart_0n );
  EO I16_I11_I5 ( I16_addOut_0n_2_, I16_I11_ha, I16_c_0n_2_ );
  EO I16_I11_I4 ( I16_I11_ha, I16_n_0n[2], z_0d[2] );
  NR2 I16_I11_I1 ( I16_I11_cv, I16_nStart_0n, I16_nCv_0n_2_ );
  IV I16_I11_I0 ( I16_I11_start, I16_nStart_0n );
  EO I16_I12_I5 ( I16_addOut_0n_3_, I16_I12_ha, I16_c_0n_3_ );
  EO I16_I12_I4 ( I16_I12_ha, I16_n_0n[3], z_0d[3] );
  NR2 I16_I12_I1 ( I16_I12_cv, I16_nStart_0n, I16_nCv_0n_3_ );
  IV I16_I12_I0 ( I16_I12_start, I16_nStart_0n );
  EO I16_I13_I5 ( I16_addOut_0n_4_, I16_I13_ha, I16_c_0n_4_ );
  EO I16_I13_I4 ( I16_I13_ha, I16_n_0n[4], z_0d[4] );
  NR2 I16_I13_I1 ( I16_I13_cv, I16_nStart_0n, I16_nCv_0n_4_ );
  IV I16_I13_I0 ( I16_I13_start, I16_nStart_0n );
  EO I16_I14_I5 ( I16_addOut_0n_5_, I16_I14_ha, I16_c_0n_5_ );
  EO I16_I14_I4 ( I16_I14_ha, I16_n_0n[5], z_0d[5] );
  NR2 I16_I14_I1 ( I16_I14_cv, I16_nStart_0n, I16_nCv_0n_5_ );
  IV I16_I14_I0 ( I16_I14_start, I16_nStart_0n );
  EO I16_I15_I5 ( I16_addOut_0n_6_, I16_I15_ha, I16_c_0n_6_ );
  EO I16_I15_I4 ( I16_I15_ha, I16_n_0n[6], z_0d[6] );
  NR2 I16_I15_I1 ( I16_I15_cv, I16_nStart_0n, I16_nCv_0n_6_ );
  IV I16_I15_I0 ( I16_I15_start, I16_nStart_0n );
  EO I16_I16_I5 ( I16_addOut_0n_7_, I16_I16_ha, I16_c_0n_7_ );
  EO I16_I16_I4 ( I16_I16_ha, I16_n_0n[7], z_0d[7] );
  NR2 I16_I16_I1 ( I16_I16_cv, I16_nStart_0n, I16_nCv_0n_7_ );
  IV I16_I16_I0 ( I16_I16_start, I16_nStart_0n );
  EO I21_I11_I5 ( c18_d[0], I21_I11_ha, I21_vcc );
  EO I21_I11_I4 ( I21_I11_ha, I21_n_0n[0], z_0d[0] );
  NR2 I21_I11_I1 ( I21_I11_cv, I21_nStart_0n, I21_nStart_0n );
  IV I21_I11_I0 ( I21_I11_start, I21_nStart_0n );
  EO I21_I12_I5 ( c18_d[1], I21_I12_ha, I21_c_0n[1] );
  EO I21_I12_I4 ( I21_I12_ha, I21_n_0n[1], z_0d[1] );
  NR2 I21_I12_I1 ( I21_I12_cv, I21_nStart_0n, I21_nCv_0n_1_ );
  IV I21_I12_I0 ( I21_I12_start, I21_nStart_0n );
  EO I21_I13_I5 ( c18_d[2], I21_I13_ha, I21_c_0n[2] );
  EO I21_I13_I4 ( I21_I13_ha, I21_n_0n[2], z_0d[2] );
  NR2 I21_I13_I1 ( I21_I13_cv, I21_nStart_0n, I21_nCv_0n_2_ );
  IV I21_I13_I0 ( I21_I13_start, I21_nStart_0n );
  EO I21_I14_I5 ( c18_d[3], I21_I14_ha, I21_c_0n[3] );
  EO I21_I14_I4 ( I21_I14_ha, I21_n_0n[3], z_0d[3] );
  NR2 I21_I14_I1 ( I21_I14_cv, I21_nStart_0n, I21_nCv_0n_3_ );
  IV I21_I14_I0 ( I21_I14_start, I21_nStart_0n );
  EO I21_I15_I5 ( c18_d[4], I21_I15_ha, I21_c_0n[4] );
  EO I21_I15_I4 ( I21_I15_ha, I21_n_0n[4], z_0d[4] );
  NR2 I21_I15_I1 ( I21_I15_cv, I21_nStart_0n, I21_nCv_0n_4_ );
  IV I21_I15_I0 ( I21_I15_start, I21_nStart_0n );
  EO I21_I16_I5 ( c18_d[5], I21_I16_ha, I21_c_0n[5] );
  EO I21_I16_I4 ( I21_I16_ha, I21_n_0n[5], z_0d[5] );
  NR2 I21_I16_I1 ( I21_I16_cv, I21_nStart_0n, I21_nCv_0n_5_ );
  IV I21_I16_I0 ( I21_I16_start, I21_nStart_0n );
  EO I21_I17_I5 ( c18_d[6], I21_I17_ha, I21_c_0n[6] );
  EO I21_I17_I4 ( I21_I17_ha, I21_n_0n[6], z_0d[6] );
  NR2 I21_I17_I1 ( I21_I17_cv, I21_nStart_0n, I21_nCv_0n_6_ );
  IV I21_I17_I0 ( I21_I17_start, I21_nStart_0n );
  EO I21_I18_I5 ( c18_d[7], I21_I18_ha, I21_c_0n[7] );
  EO I21_I18_I4 ( I21_I18_ha, I21_n_0n[7], z_0d[7] );
  NR2 I21_I18_I1 ( I21_I18_cv, I21_nStart_0n, I21_nCv_0n_7_ );
  IV I21_I18_I0 ( I21_I18_start, I21_nStart_0n );
  EO I26_I11_I5 ( c9_d[0], I26_I11_ha, I26_vcc );
  EO I26_I11_I4 ( I26_I11_ha, I26_n_0n[0], c34_d[0] );
  NR2 I26_I11_I1 ( I26_I11_cv, I26_nStart_0n, I26_nStart_0n );
  IV I26_I11_I0 ( I26_I11_start, I26_nStart_0n );
  EO I26_I12_I5 ( c9_d[1], I26_I12_ha, I26_c_0n[1] );
  EO I26_I12_I4 ( I26_I12_ha, I26_n_0n[1], c34_d[1] );
  NR2 I26_I12_I1 ( I26_I12_cv, I26_nStart_0n, I26_nCv_0n_1_ );
  IV I26_I12_I0 ( I26_I12_start, I26_nStart_0n );
  EO I26_I13_I5 ( c9_d[2], I26_I13_ha, I26_c_0n[2] );
  EO I26_I13_I4 ( I26_I13_ha, I26_n_0n[2], c34_d[2] );
  NR2 I26_I13_I1 ( I26_I13_cv, I26_nStart_0n, I26_nCv_0n_2_ );
  IV I26_I13_I0 ( I26_I13_start, I26_nStart_0n );
  EO I26_I14_I5 ( c9_d[3], I26_I14_ha, I26_c_0n[3] );
  EO I26_I14_I4 ( I26_I14_ha, I26_n_0n[3], c34_d[3] );
  NR2 I26_I14_I1 ( I26_I14_cv, I26_nStart_0n, I26_nCv_0n_3_ );
  IV I26_I14_I0 ( I26_I14_start, I26_nStart_0n );
  EO I26_I15_I5 ( c9_d[4], I26_I15_ha, I26_c_0n[4] );
  EO I26_I15_I4 ( I26_I15_ha, I26_n_0n[4], c34_d[4] );
  NR2 I26_I15_I1 ( I26_I15_cv, I26_nStart_0n, I26_nCv_0n_4_ );
  IV I26_I15_I0 ( I26_I15_start, I26_nStart_0n );
  EO I26_I16_I5 ( c9_d[5], I26_I16_ha, I26_c_0n[5] );
  EO I26_I16_I4 ( I26_I16_ha, I26_n_0n[5], c34_d[5] );
  NR2 I26_I16_I1 ( I26_I16_cv, I26_nStart_0n, I26_nCv_0n_5_ );
  IV I26_I16_I0 ( I26_I16_start, I26_nStart_0n );
  EO I26_I17_I5 ( c9_d[6], I26_I17_ha, I26_c_0n[6] );
  EO I26_I17_I4 ( I26_I17_ha, I26_n_0n[6], c34_d[6] );
  NR2 I26_I17_I1 ( I26_I17_cv, I26_nStart_0n, I26_nCv_0n_6_ );
  IV I26_I17_I0 ( I26_I17_start, I26_nStart_0n );
  EO I26_I18_I5 ( c9_d[7], I26_I18_ha, I26_c_0n[7] );
  EO I26_I18_I4 ( I26_I18_ha, I26_n_0n[7], c34_d[7] );
  NR2 I26_I18_I1 ( I26_I18_cv, I26_nStart_0n, I26_nCv_0n_7_ );
  IV I26_I18_I0 ( I26_I18_start, I26_nStart_0n );
  IV I16_I9_I2_I1 ( I16_I9_I2_nsel_0n, I16_I9_ha );
  IV I16_I10_I2_I1 ( I16_I10_I2_nsel_0n, I16_I10_ha );
  IV I16_I11_I2_I1 ( I16_I11_I2_nsel_0n, I16_I11_ha );
  IV I16_I12_I2_I1 ( I16_I12_I2_nsel_0n, I16_I12_ha );
  IV I16_I13_I2_I1 ( I16_I13_I2_nsel_0n, I16_I13_ha );
  IV I16_I14_I2_I1 ( I16_I14_I2_nsel_0n, I16_I14_ha );
  IV I16_I15_I2_I1 ( I16_I15_I2_nsel_0n, I16_I15_ha );
  IV I16_I16_I2_I1 ( I16_I16_I2_nsel_0n, I16_I16_ha );
  IV I21_I11_I2_I1 ( I21_I11_I2_nsel_0n, I21_I11_ha );
  IV I21_I12_I2_I1 ( I21_I12_I2_nsel_0n, I21_I12_ha );
  IV I21_I13_I2_I1 ( I21_I13_I2_nsel_0n, I21_I13_ha );
  IV I21_I14_I2_I1 ( I21_I14_I2_nsel_0n, I21_I14_ha );
  IV I21_I15_I2_I1 ( I21_I15_I2_nsel_0n, I21_I15_ha );
  IV I21_I16_I2_I1 ( I21_I16_I2_nsel_0n, I21_I16_ha );
  IV I21_I17_I2_I1 ( I21_I17_I2_nsel_0n, I21_I17_ha );
  IV I21_I18_I2_I1 ( I21_I18_I2_nsel_0n, I21_I18_ha );
  IV I26_I11_I2_I1 ( I26_I11_I2_nsel_0n, I26_I11_ha );
  IV I26_I12_I2_I1 ( I26_I12_I2_nsel_0n, I26_I12_ha );
  IV I26_I13_I2_I1 ( I26_I13_I2_nsel_0n, I26_I13_ha );
  IV I26_I14_I2_I1 ( I26_I14_I2_nsel_0n, I26_I14_ha );
  IV I26_I15_I2_I1 ( I26_I15_I2_nsel_0n, I26_I15_ha );
  IV I26_I16_I2_I1 ( I26_I16_I2_nsel_0n, I26_I16_ha );
  IV I26_I17_I2_I1 ( I26_I17_I2_nsel_0n, I26_I17_ha );
  IV I26_I18_I2_I1 ( I26_I18_I2_nsel_0n, I26_I18_ha );
  AN2 I16_I9_I2_I0_I2 ( I16_I9_I2_I0_int_0n[0], I16_I9_start, I16_I9_I2_nsel_0n );
  AN2 I16_I9_I2_I0_I1 ( I16_I9_I2_I0_int_0n[1], I16_I9_cv, I16_I9_ha );
  NR2 I16_I9_I2_I0_I0 ( I16_nCv_0n_1_, I16_I9_I2_I0_int_0n[0], I16_I9_I2_I0_int_0n[1] );
  AN2 I16_I10_I2_I0_I2 ( I16_I10_I2_I0_int_0n[0], I16_I10_start, I16_I10_I2_nsel_0n );
  AN2 I16_I10_I2_I0_I1 ( I16_I10_I2_I0_int_0n[1], I16_I10_cv, I16_I10_ha );
  NR2 I16_I10_I2_I0_I0 ( I16_nCv_0n_2_, I16_I10_I2_I0_int_0n[0], I16_I10_I2_I0_int_0n[1] );
  AN2 I16_I11_I2_I0_I2 ( I16_I11_I2_I0_int_0n[0], I16_I11_start, I16_I11_I2_nsel_0n );
  AN2 I16_I11_I2_I0_I1 ( I16_I11_I2_I0_int_0n[1], I16_I11_cv, I16_I11_ha );
  NR2 I16_I11_I2_I0_I0 ( I16_nCv_0n_3_, I16_I11_I2_I0_int_0n[0], I16_I11_I2_I0_int_0n[1] );
  AN2 I16_I12_I2_I0_I2 ( I16_I12_I2_I0_int_0n[0], I16_I12_start, I16_I12_I2_nsel_0n );
  AN2 I16_I12_I2_I0_I1 ( I16_I12_I2_I0_int_0n[1], I16_I12_cv, I16_I12_ha );
  NR2 I16_I12_I2_I0_I0 ( I16_nCv_0n_4_, I16_I12_I2_I0_int_0n[0], I16_I12_I2_I0_int_0n[1] );
  AN2 I16_I13_I2_I0_I2 ( I16_I13_I2_I0_int_0n[0], I16_I13_start, I16_I13_I2_nsel_0n );
  AN2 I16_I13_I2_I0_I1 ( I16_I13_I2_I0_int_0n[1], I16_I13_cv, I16_I13_ha );
  NR2 I16_I13_I2_I0_I0 ( I16_nCv_0n_5_, I16_I13_I2_I0_int_0n[0], I16_I13_I2_I0_int_0n[1] );
  AN2 I16_I14_I2_I0_I2 ( I16_I14_I2_I0_int_0n[0], I16_I14_start, I16_I14_I2_nsel_0n );
  AN2 I16_I14_I2_I0_I1 ( I16_I14_I2_I0_int_0n[1], I16_I14_cv, I16_I14_ha );
  NR2 I16_I14_I2_I0_I0 ( I16_nCv_0n_6_, I16_I14_I2_I0_int_0n[0], I16_I14_I2_I0_int_0n[1] );
  AN2 I16_I15_I2_I0_I2 ( I16_I15_I2_I0_int_0n[0], I16_I15_start, I16_I15_I2_nsel_0n );
  AN2 I16_I15_I2_I0_I1 ( I16_I15_I2_I0_int_0n[1], I16_I15_cv, I16_I15_ha );
  NR2 I16_I15_I2_I0_I0 ( I16_nCv_0n_7_, I16_I15_I2_I0_int_0n[0], I16_I15_I2_I0_int_0n[1] );
  AN2 I16_I16_I2_I0_I2 ( I16_I16_I2_I0_int_0n[0], I16_I16_start, I16_I16_I2_nsel_0n );
  AN2 I16_I16_I2_I0_I1 ( I16_I16_I2_I0_int_0n[1], I16_I16_cv, I16_I16_ha );
  NR2 I16_I16_I2_I0_I0 ( I16_nCv_0n_8_, I16_I16_I2_I0_int_0n[0], I16_I16_I2_I0_int_0n[1] );
  AN2 I21_I11_I2_I0_I2 ( I21_I11_I2_I0_int_0n[0], I21_I11_start, I21_I11_I2_nsel_0n );
  AN2 I21_I11_I2_I0_I1 ( I21_I11_I2_I0_int_0n[1], I21_I11_cv, I21_I11_ha );
  NR2 I21_I11_I2_I0_I0 ( I21_nCv_0n_1_, I21_I11_I2_I0_int_0n[0], I21_I11_I2_I0_int_0n[1] );
  AN2 I21_I12_I2_I0_I2 ( I21_I12_I2_I0_int_0n[0], I21_I12_start, I21_I12_I2_nsel_0n );
  AN2 I21_I12_I2_I0_I1 ( I21_I12_I2_I0_int_0n[1], I21_I12_cv, I21_I12_ha );
  NR2 I21_I12_I2_I0_I0 ( I21_nCv_0n_2_, I21_I12_I2_I0_int_0n[0], I21_I12_I2_I0_int_0n[1] );
  AN2 I21_I13_I2_I0_I2 ( I21_I13_I2_I0_int_0n[0], I21_I13_start, I21_I13_I2_nsel_0n );
  AN2 I21_I13_I2_I0_I1 ( I21_I13_I2_I0_int_0n[1], I21_I13_cv, I21_I13_ha );
  NR2 I21_I13_I2_I0_I0 ( I21_nCv_0n_3_, I21_I13_I2_I0_int_0n[0], I21_I13_I2_I0_int_0n[1] );
  AN2 I21_I14_I2_I0_I2 ( I21_I14_I2_I0_int_0n[0], I21_I14_start, I21_I14_I2_nsel_0n );
  AN2 I21_I14_I2_I0_I1 ( I21_I14_I2_I0_int_0n[1], I21_I14_cv, I21_I14_ha );
  NR2 I21_I14_I2_I0_I0 ( I21_nCv_0n_4_, I21_I14_I2_I0_int_0n[0], I21_I14_I2_I0_int_0n[1] );
  AN2 I21_I15_I2_I0_I2 ( I21_I15_I2_I0_int_0n[0], I21_I15_start, I21_I15_I2_nsel_0n );
  AN2 I21_I15_I2_I0_I1 ( I21_I15_I2_I0_int_0n[1], I21_I15_cv, I21_I15_ha );
  NR2 I21_I15_I2_I0_I0 ( I21_nCv_0n_5_, I21_I15_I2_I0_int_0n[0], I21_I15_I2_I0_int_0n[1] );
  AN2 I21_I16_I2_I0_I2 ( I21_I16_I2_I0_int_0n[0], I21_I16_start, I21_I16_I2_nsel_0n );
  AN2 I21_I16_I2_I0_I1 ( I21_I16_I2_I0_int_0n[1], I21_I16_cv, I21_I16_ha );
  NR2 I21_I16_I2_I0_I0 ( I21_nCv_0n_6_, I21_I16_I2_I0_int_0n[0], I21_I16_I2_I0_int_0n[1] );
  AN2 I21_I17_I2_I0_I2 ( I21_I17_I2_I0_int_0n[0], I21_I17_start, I21_I17_I2_nsel_0n );
  AN2 I21_I17_I2_I0_I1 ( I21_I17_I2_I0_int_0n[1], I21_I17_cv, I21_I17_ha );
  NR2 I21_I17_I2_I0_I0 ( I21_nCv_0n_7_, I21_I17_I2_I0_int_0n[0], I21_I17_I2_I0_int_0n[1] );
  AN2 I21_I18_I2_I0_I2 ( I21_I18_I2_I0_int_0n[0], I21_I18_start, I21_I18_I2_nsel_0n );
  AN2 I21_I18_I2_I0_I1 ( I21_I18_I2_I0_int_0n[1], I21_I18_cv, I21_I18_ha );
  NR2 I21_I18_I2_I0_I0 ( I21_nCv_0n_8_, I21_I18_I2_I0_int_0n[0], I21_I18_I2_I0_int_0n[1] );
  AN2 I26_I11_I2_I0_I2 ( I26_I11_I2_I0_int_0n[0], I26_I11_start, I26_I11_I2_nsel_0n );
  AN2 I26_I11_I2_I0_I1 ( I26_I11_I2_I0_int_0n[1], I26_I11_cv, I26_I11_ha );
  NR2 I26_I11_I2_I0_I0 ( I26_nCv_0n_1_, I26_I11_I2_I0_int_0n[0], I26_I11_I2_I0_int_0n[1] );
  AN2 I26_I12_I2_I0_I2 ( I26_I12_I2_I0_int_0n[0], I26_I12_start, I26_I12_I2_nsel_0n );
  AN2 I26_I12_I2_I0_I1 ( I26_I12_I2_I0_int_0n[1], I26_I12_cv, I26_I12_ha );
  NR2 I26_I12_I2_I0_I0 ( I26_nCv_0n_2_, I26_I12_I2_I0_int_0n[0], I26_I12_I2_I0_int_0n[1] );
  AN2 I26_I13_I2_I0_I2 ( I26_I13_I2_I0_int_0n[0], I26_I13_start, I26_I13_I2_nsel_0n );
  AN2 I26_I13_I2_I0_I1 ( I26_I13_I2_I0_int_0n[1], I26_I13_cv, I26_I13_ha );
  NR2 I26_I13_I2_I0_I0 ( I26_nCv_0n_3_, I26_I13_I2_I0_int_0n[0], I26_I13_I2_I0_int_0n[1] );
  AN2 I26_I14_I2_I0_I2 ( I26_I14_I2_I0_int_0n[0], I26_I14_start, I26_I14_I2_nsel_0n );
  AN2 I26_I14_I2_I0_I1 ( I26_I14_I2_I0_int_0n[1], I26_I14_cv, I26_I14_ha );
  NR2 I26_I14_I2_I0_I0 ( I26_nCv_0n_4_, I26_I14_I2_I0_int_0n[0], I26_I14_I2_I0_int_0n[1] );
  AN2 I26_I15_I2_I0_I2 ( I26_I15_I2_I0_int_0n[0], I26_I15_start, I26_I15_I2_nsel_0n );
  AN2 I26_I15_I2_I0_I1 ( I26_I15_I2_I0_int_0n[1], I26_I15_cv, I26_I15_ha );
  NR2 I26_I15_I2_I0_I0 ( I26_nCv_0n_5_, I26_I15_I2_I0_int_0n[0], I26_I15_I2_I0_int_0n[1] );
  AN2 I26_I16_I2_I0_I2 ( I26_I16_I2_I0_int_0n[0], I26_I16_start, I26_I16_I2_nsel_0n );
  AN2 I26_I16_I2_I0_I1 ( I26_I16_I2_I0_int_0n[1], I26_I16_cv, I26_I16_ha );
  NR2 I26_I16_I2_I0_I0 ( I26_nCv_0n_6_, I26_I16_I2_I0_int_0n[0], I26_I16_I2_I0_int_0n[1] );
  AN2 I26_I17_I2_I0_I2 ( I26_I17_I2_I0_int_0n[0], I26_I17_start, I26_I17_I2_nsel_0n );
  AN2 I26_I17_I2_I0_I1 ( I26_I17_I2_I0_int_0n[1], I26_I17_cv, I26_I17_ha );
  NR2 I26_I17_I2_I0_I0 ( I26_nCv_0n_7_, I26_I17_I2_I0_int_0n[0], I26_I17_I2_I0_int_0n[1] );
  AN2 I26_I18_I2_I0_I2 ( I26_I18_I2_I0_int_0n[0], I26_I18_start, I26_I18_I2_nsel_0n );
  AN2 I26_I18_I2_I0_I1 ( I26_I18_I2_I0_int_0n[1], I26_I18_cv, I26_I18_ha );
  NR2 I26_I18_I2_I0_I0 ( I26_nCv_0n_8_, I26_I18_I2_I0_int_0n[0], I26_I18_I2_I0_int_0n[1] );
  IV I1_I0_I1 ( I1_I0_nsel_0n, I1_select_0n );
  IV I1_I1_I1 ( I1_I1_nsel_0n, I1_select_0n );
  IV I1_I2_I1 ( I1_I2_nsel_0n, I1_select_0n );
  IV I1_I3_I1 ( I1_I3_nsel_0n, I1_select_0n );
  IV I1_I4_I1 ( I1_I4_nsel_0n, I1_select_0n );
  IV I1_I5_I1 ( I1_I5_nsel_0n, I1_select_0n );
  IV I1_I6_I1 ( I1_I6_nsel_0n, I1_select_0n );
  IV I1_I7_I1 ( I1_I7_nsel_0n, I1_select_0n );
  IV I1_I8_I1 ( I1_I8_nsel_0n, I1_select_0n );
  IV I3_I0_I1 ( I3_I0_nsel_0n, I3_select_0n );
  IV I3_I1_I1 ( I3_I1_nsel_0n, I3_select_0n );
  IV I3_I2_I1 ( I3_I2_nsel_0n, I3_select_0n );
  IV I3_I3_I1 ( I3_I3_nsel_0n, I3_select_0n );
  IV I3_I4_I1 ( I3_I4_nsel_0n, I3_select_0n );
  IV I3_I5_I1 ( I3_I5_nsel_0n, I3_select_0n );
  IV I3_I6_I1 ( I3_I6_nsel_0n, I3_select_0n );
  IV I3_I7_I1 ( I3_I7_nsel_0n, I3_select_0n );
  IV I3_I8_I1 ( I3_I8_nsel_0n, I3_select_0n );
  IV I16_I9_I3_I1 ( I16_I9_I3_nsel_0n, I16_I9_ha );
  IV I16_I10_I3_I1 ( I16_I10_I3_nsel_0n, I16_I10_ha );
  IV I16_I11_I3_I1 ( I16_I11_I3_nsel_0n, I16_I11_ha );
  IV I16_I12_I3_I1 ( I16_I12_I3_nsel_0n, I16_I12_ha );
  IV I16_I13_I3_I1 ( I16_I13_I3_nsel_0n, I16_I13_ha );
  IV I16_I14_I3_I1 ( I16_I14_I3_nsel_0n, I16_I14_ha );
  IV I16_I15_I3_I1 ( I16_I15_I3_nsel_0n, I16_I15_ha );
  IV I16_I16_I3_I1 ( I16_I16_I3_nsel_0n, I16_I16_ha );
  IV I21_I11_I3_I1 ( I21_I11_I3_nsel_0n, I21_I11_ha );
  IV I21_I12_I3_I1 ( I21_I12_I3_nsel_0n, I21_I12_ha );
  IV I21_I13_I3_I1 ( I21_I13_I3_nsel_0n, I21_I13_ha );
  IV I21_I14_I3_I1 ( I21_I14_I3_nsel_0n, I21_I14_ha );
  IV I21_I15_I3_I1 ( I21_I15_I3_nsel_0n, I21_I15_ha );
  IV I21_I16_I3_I1 ( I21_I16_I3_nsel_0n, I21_I16_ha );
  IV I21_I17_I3_I1 ( I21_I17_I3_nsel_0n, I21_I17_ha );
  IV I21_I18_I3_I1 ( I21_I18_I3_nsel_0n, I21_I18_ha );
  IV I26_I11_I3_I1 ( I26_I11_I3_nsel_0n, I26_I11_ha );
  IV I26_I12_I3_I1 ( I26_I12_I3_nsel_0n, I26_I12_ha );
  IV I26_I13_I3_I1 ( I26_I13_I3_nsel_0n, I26_I13_ha );
  IV I26_I14_I3_I1 ( I26_I14_I3_nsel_0n, I26_I14_ha );
  IV I26_I15_I3_I1 ( I26_I15_I3_nsel_0n, I26_I15_ha );
  IV I26_I16_I3_I1 ( I26_I16_I3_nsel_0n, I26_I16_ha );
  IV I26_I17_I3_I1 ( I26_I17_I3_nsel_0n, I26_I17_ha );
  IV I26_I18_I3_I1 ( I26_I18_I3_nsel_0n, I26_I18_ha );
  AN2 I1_I0_I0_I2 ( I1_I0_I0_int_0n[0], c24_d[0], I1_I0_nsel_0n );
  AN2 I1_I0_I0_I1 ( I1_I0_I0_int_0n[1], x_0d[0], I1_select_0n );
  OR2 I1_I0_I0_I0 ( c45_d[0], I1_I0_I0_int_0n[0], I1_I0_I0_int_0n[1] );
  AN2 I1_I1_I0_I2 ( I1_I1_I0_int_0n[0], c24_d[1], I1_I1_nsel_0n );
  AN2 I1_I1_I0_I1 ( I1_I1_I0_int_0n[1], x_0d[1], I1_select_0n );
  OR2 I1_I1_I0_I0 ( c45_d[1], I1_I1_I0_int_0n[0], I1_I1_I0_int_0n[1] );
  AN2 I1_I2_I0_I2 ( I1_I2_I0_int_0n[0], c24_d[2], I1_I2_nsel_0n );
  AN2 I1_I2_I0_I1 ( I1_I2_I0_int_0n[1], x_0d[2], I1_select_0n );
  OR2 I1_I2_I0_I0 ( c45_d[2], I1_I2_I0_int_0n[0], I1_I2_I0_int_0n[1] );
  AN2 I1_I3_I0_I2 ( I1_I3_I0_int_0n[0], c24_d[3], I1_I3_nsel_0n );
  AN2 I1_I3_I0_I1 ( I1_I3_I0_int_0n[1], x_0d[3], I1_select_0n );
  OR2 I1_I3_I0_I0 ( c45_d[3], I1_I3_I0_int_0n[0], I1_I3_I0_int_0n[1] );
  AN2 I1_I4_I0_I2 ( I1_I4_I0_int_0n[0], c24_d[4], I1_I4_nsel_0n );
  AN2 I1_I4_I0_I1 ( I1_I4_I0_int_0n[1], x_0d[4], I1_select_0n );
  OR2 I1_I4_I0_I0 ( c45_d[4], I1_I4_I0_int_0n[0], I1_I4_I0_int_0n[1] );
  AN2 I1_I5_I0_I2 ( I1_I5_I0_int_0n[0], c24_d[5], I1_I5_nsel_0n );
  AN2 I1_I5_I0_I1 ( I1_I5_I0_int_0n[1], x_0d[5], I1_select_0n );
  OR2 I1_I5_I0_I0 ( c45_d[5], I1_I5_I0_int_0n[0], I1_I5_I0_int_0n[1] );
  AN2 I1_I6_I0_I2 ( I1_I6_I0_int_0n[0], c24_d[6], I1_I6_nsel_0n );
  AN2 I1_I6_I0_I1 ( I1_I6_I0_int_0n[1], x_0d[6], I1_select_0n );
  OR2 I1_I6_I0_I0 ( c45_d[6], I1_I6_I0_int_0n[0], I1_I6_I0_int_0n[1] );
  AN2 I1_I7_I0_I2 ( I1_I7_I0_int_0n[0], c24_d[7], I1_I7_nsel_0n );
  AN2 I1_I7_I0_I1 ( I1_I7_I0_int_0n[1], x_0d[7], I1_select_0n );
  OR2 I1_I7_I0_I0 ( c45_d[7], I1_I7_I0_int_0n[0], I1_I7_I0_int_0n[1] );
  AN2 I1_I8_I0_I2 ( I1_I8_I0_int_0n[0], c22_r, I1_I8_nsel_0n );
  AN2 I1_I8_I0_I1 ( I1_I8_I0_int_0n[1], x_0a, I1_select_0n );
  OR2 I1_I8_I0_I0 ( c45_r, I1_I8_I0_int_0n[0], I1_I8_I0_int_0n[1] );
  AN2 I3_I0_I0_I2 ( I3_I0_I0_int_0n[0], c15_d[0], I3_I0_nsel_0n );
  AN2 I3_I0_I0_I1 ( I3_I0_I0_int_0n[1], y_0d[0], I3_select_0n );
  OR2 I3_I0_I0_I0 ( c44_d[0], I3_I0_I0_int_0n[0], I3_I0_I0_int_0n[1] );
  AN2 I3_I1_I0_I2 ( I3_I1_I0_int_0n[0], c15_d[1], I3_I1_nsel_0n );
  AN2 I3_I1_I0_I1 ( I3_I1_I0_int_0n[1], y_0d[1], I3_select_0n );
  OR2 I3_I1_I0_I0 ( c44_d[1], I3_I1_I0_int_0n[0], I3_I1_I0_int_0n[1] );
  AN2 I3_I2_I0_I2 ( I3_I2_I0_int_0n[0], c15_d[2], I3_I2_nsel_0n );
  AN2 I3_I2_I0_I1 ( I3_I2_I0_int_0n[1], y_0d[2], I3_select_0n );
  OR2 I3_I2_I0_I0 ( c44_d[2], I3_I2_I0_int_0n[0], I3_I2_I0_int_0n[1] );
  AN2 I3_I3_I0_I2 ( I3_I3_I0_int_0n[0], c15_d[3], I3_I3_nsel_0n );
  AN2 I3_I3_I0_I1 ( I3_I3_I0_int_0n[1], y_0d[3], I3_select_0n );
  OR2 I3_I3_I0_I0 ( c44_d[3], I3_I3_I0_int_0n[0], I3_I3_I0_int_0n[1] );
  AN2 I3_I4_I0_I2 ( I3_I4_I0_int_0n[0], c15_d[4], I3_I4_nsel_0n );
  AN2 I3_I4_I0_I1 ( I3_I4_I0_int_0n[1], y_0d[4], I3_select_0n );
  OR2 I3_I4_I0_I0 ( c44_d[4], I3_I4_I0_int_0n[0], I3_I4_I0_int_0n[1] );
  AN2 I3_I5_I0_I2 ( I3_I5_I0_int_0n[0], c15_d[5], I3_I5_nsel_0n );
  AN2 I3_I5_I0_I1 ( I3_I5_I0_int_0n[1], y_0d[5], I3_select_0n );
  OR2 I3_I5_I0_I0 ( c44_d[5], I3_I5_I0_int_0n[0], I3_I5_I0_int_0n[1] );
  AN2 I3_I6_I0_I2 ( I3_I6_I0_int_0n[0], c15_d[6], I3_I6_nsel_0n );
  AN2 I3_I6_I0_I1 ( I3_I6_I0_int_0n[1], y_0d[6], I3_select_0n );
  OR2 I3_I6_I0_I0 ( c44_d[6], I3_I6_I0_int_0n[0], I3_I6_I0_int_0n[1] );
  AN2 I3_I7_I0_I2 ( I3_I7_I0_int_0n[0], c15_d[7], I3_I7_nsel_0n );
  AN2 I3_I7_I0_I1 ( I3_I7_I0_int_0n[1], y_0d[7], I3_select_0n );
  OR2 I3_I7_I0_I0 ( c44_d[7], I3_I7_I0_int_0n[0], I3_I7_I0_int_0n[1] );
  AN2 I3_I8_I0_I2 ( I3_I8_I0_int_0n[0], c13_r, I3_I8_nsel_0n );
  AN2 I3_I8_I0_I1 ( I3_I8_I0_int_0n[1], y_0a, I3_select_0n );
  OR2 I3_I8_I0_I0 ( c44_r, I3_I8_I0_int_0n[0], I3_I8_I0_int_0n[1] );
  AN2 I16_I9_I3_I0_I2 ( I16_I9_I3_I0_int_0n[0], I16_n_0n[0], I16_I9_I3_nsel_0n );
  AN2 I16_I9_I3_I0_I1 ( I16_I9_I3_I0_int_0n[1], I16_vcc, I16_I9_ha );
  OR2 I16_I9_I3_I0_I0 ( I16_c_0n_1_, I16_I9_I3_I0_int_0n[0], I16_I9_I3_I0_int_0n[1] );
  AN2 I16_I10_I3_I0_I2 ( I16_I10_I3_I0_int_0n[0], I16_n_0n[1], I16_I10_I3_nsel_0n );
  AN2 I16_I10_I3_I0_I1 ( I16_I10_I3_I0_int_0n[1], I16_c_0n_1_, I16_I10_ha );
  OR2 I16_I10_I3_I0_I0 ( I16_c_0n_2_, I16_I10_I3_I0_int_0n[0], I16_I10_I3_I0_int_0n[1] );
  AN2 I16_I11_I3_I0_I2 ( I16_I11_I3_I0_int_0n[0], I16_n_0n[2], I16_I11_I3_nsel_0n );
  AN2 I16_I11_I3_I0_I1 ( I16_I11_I3_I0_int_0n[1], I16_c_0n_2_, I16_I11_ha );
  OR2 I16_I11_I3_I0_I0 ( I16_c_0n_3_, I16_I11_I3_I0_int_0n[0], I16_I11_I3_I0_int_0n[1] );
  AN2 I16_I12_I3_I0_I2 ( I16_I12_I3_I0_int_0n[0], I16_n_0n[3], I16_I12_I3_nsel_0n );
  AN2 I16_I12_I3_I0_I1 ( I16_I12_I3_I0_int_0n[1], I16_c_0n_3_, I16_I12_ha );
  OR2 I16_I12_I3_I0_I0 ( I16_c_0n_4_, I16_I12_I3_I0_int_0n[0], I16_I12_I3_I0_int_0n[1] );
  AN2 I16_I13_I3_I0_I2 ( I16_I13_I3_I0_int_0n[0], I16_n_0n[4], I16_I13_I3_nsel_0n );
  AN2 I16_I13_I3_I0_I1 ( I16_I13_I3_I0_int_0n[1], I16_c_0n_4_, I16_I13_ha );
  OR2 I16_I13_I3_I0_I0 ( I16_c_0n_5_, I16_I13_I3_I0_int_0n[0], I16_I13_I3_I0_int_0n[1] );
  AN2 I16_I14_I3_I0_I2 ( I16_I14_I3_I0_int_0n[0], I16_n_0n[5], I16_I14_I3_nsel_0n );
  AN2 I16_I14_I3_I0_I1 ( I16_I14_I3_I0_int_0n[1], I16_c_0n_5_, I16_I14_ha );
  OR2 I16_I14_I3_I0_I0 ( I16_c_0n_6_, I16_I14_I3_I0_int_0n[0], I16_I14_I3_I0_int_0n[1] );
  AN2 I16_I15_I3_I0_I2 ( I16_I15_I3_I0_int_0n[0], I16_n_0n[6], I16_I15_I3_nsel_0n );
  AN2 I16_I15_I3_I0_I1 ( I16_I15_I3_I0_int_0n[1], I16_c_0n_6_, I16_I15_ha );
  OR2 I16_I15_I3_I0_I0 ( I16_c_0n_7_, I16_I15_I3_I0_int_0n[0], I16_I15_I3_I0_int_0n[1] );
  AN2 I16_I16_I3_I0_I2 ( I16_I16_I3_I0_int_0n[0], I16_n_0n[7], I16_I16_I3_nsel_0n );
  AN2 I16_I16_I3_I0_I1 ( I16_I16_I3_I0_int_0n[1], I16_c_0n_7_, I16_I16_ha );
  OR2 I16_I16_I3_I0_I0 ( I16_c_0n_8_, I16_I16_I3_I0_int_0n[0], I16_I16_I3_I0_int_0n[1] );
  AN2 I21_I11_I3_I0_I2 ( I21_I11_I3_I0_int_0n[0], I21_n_0n[0], I21_I11_I3_nsel_0n );
  AN2 I21_I11_I3_I0_I1 ( I21_I11_I3_I0_int_0n[1], I21_vcc, I21_I11_ha );
  OR2 I21_I11_I3_I0_I0 ( I21_c_0n[1], I21_I11_I3_I0_int_0n[0], I21_I11_I3_I0_int_0n[1] );
  AN2 I21_I12_I3_I0_I2 ( I21_I12_I3_I0_int_0n[0], I21_n_0n[1], I21_I12_I3_nsel_0n );
  AN2 I21_I12_I3_I0_I1 ( I21_I12_I3_I0_int_0n[1], I21_c_0n[1], I21_I12_ha );
  OR2 I21_I12_I3_I0_I0 ( I21_c_0n[2], I21_I12_I3_I0_int_0n[0], I21_I12_I3_I0_int_0n[1] );
  AN2 I21_I13_I3_I0_I2 ( I21_I13_I3_I0_int_0n[0], I21_n_0n[2], I21_I13_I3_nsel_0n );
  AN2 I21_I13_I3_I0_I1 ( I21_I13_I3_I0_int_0n[1], I21_c_0n[2], I21_I13_ha );
  OR2 I21_I13_I3_I0_I0 ( I21_c_0n[3], I21_I13_I3_I0_int_0n[0], I21_I13_I3_I0_int_0n[1] );
  AN2 I21_I14_I3_I0_I2 ( I21_I14_I3_I0_int_0n[0], I21_n_0n[3], I21_I14_I3_nsel_0n );
  AN2 I21_I14_I3_I0_I1 ( I21_I14_I3_I0_int_0n[1], I21_c_0n[3], I21_I14_ha );
  OR2 I21_I14_I3_I0_I0 ( I21_c_0n[4], I21_I14_I3_I0_int_0n[0], I21_I14_I3_I0_int_0n[1] );
  AN2 I21_I15_I3_I0_I2 ( I21_I15_I3_I0_int_0n[0], I21_n_0n[4], I21_I15_I3_nsel_0n );
  AN2 I21_I15_I3_I0_I1 ( I21_I15_I3_I0_int_0n[1], I21_c_0n[4], I21_I15_ha );
  OR2 I21_I15_I3_I0_I0 ( I21_c_0n[5], I21_I15_I3_I0_int_0n[0], I21_I15_I3_I0_int_0n[1] );
  AN2 I21_I16_I3_I0_I2 ( I21_I16_I3_I0_int_0n[0], I21_n_0n[5], I21_I16_I3_nsel_0n );
  AN2 I21_I16_I3_I0_I1 ( I21_I16_I3_I0_int_0n[1], I21_c_0n[5], I21_I16_ha );
  OR2 I21_I16_I3_I0_I0 ( I21_c_0n[6], I21_I16_I3_I0_int_0n[0], I21_I16_I3_I0_int_0n[1] );
  AN2 I21_I17_I3_I0_I2 ( I21_I17_I3_I0_int_0n[0], I21_n_0n[6], I21_I17_I3_nsel_0n );
  AN2 I21_I17_I3_I0_I1 ( I21_I17_I3_I0_int_0n[1], I21_c_0n[6], I21_I17_ha );
  OR2 I21_I17_I3_I0_I0 ( I21_c_0n[7], I21_I17_I3_I0_int_0n[0], I21_I17_I3_I0_int_0n[1] );
  AN2 I21_I18_I3_I0_I2 ( I21_I18_I3_I0_int_0n[0], I21_n_0n[7], I21_I18_I3_nsel_0n );
  AN2 I21_I18_I3_I0_I1 ( I21_I18_I3_I0_int_0n[1], I21_c_0n[7], I21_I18_ha );
  OR2 I21_I18_I3_I0_I0 ( I21_c_0n[8], I21_I18_I3_I0_int_0n[0], I21_I18_I3_I0_int_0n[1] );
  AN2 I26_I11_I3_I0_I2 ( I26_I11_I3_I0_int_0n[0], I26_n_0n[0], I26_I11_I3_nsel_0n );
  AN2 I26_I11_I3_I0_I1 ( I26_I11_I3_I0_int_0n[1], I26_vcc, I26_I11_ha );
  OR2 I26_I11_I3_I0_I0 ( I26_c_0n[1], I26_I11_I3_I0_int_0n[0], I26_I11_I3_I0_int_0n[1] );
  AN2 I26_I12_I3_I0_I2 ( I26_I12_I3_I0_int_0n[0], I26_n_0n[1], I26_I12_I3_nsel_0n );
  AN2 I26_I12_I3_I0_I1 ( I26_I12_I3_I0_int_0n[1], I26_c_0n[1], I26_I12_ha );
  OR2 I26_I12_I3_I0_I0 ( I26_c_0n[2], I26_I12_I3_I0_int_0n[0], I26_I12_I3_I0_int_0n[1] );
  AN2 I26_I13_I3_I0_I2 ( I26_I13_I3_I0_int_0n[0], I26_n_0n[2], I26_I13_I3_nsel_0n );
  AN2 I26_I13_I3_I0_I1 ( I26_I13_I3_I0_int_0n[1], I26_c_0n[2], I26_I13_ha );
  OR2 I26_I13_I3_I0_I0 ( I26_c_0n[3], I26_I13_I3_I0_int_0n[0], I26_I13_I3_I0_int_0n[1] );
  AN2 I26_I14_I3_I0_I2 ( I26_I14_I3_I0_int_0n[0], I26_n_0n[3], I26_I14_I3_nsel_0n );
  AN2 I26_I14_I3_I0_I1 ( I26_I14_I3_I0_int_0n[1], I26_c_0n[3], I26_I14_ha );
  OR2 I26_I14_I3_I0_I0 ( I26_c_0n[4], I26_I14_I3_I0_int_0n[0], I26_I14_I3_I0_int_0n[1] );
  AN2 I26_I15_I3_I0_I2 ( I26_I15_I3_I0_int_0n[0], I26_n_0n[4], I26_I15_I3_nsel_0n );
  AN2 I26_I15_I3_I0_I1 ( I26_I15_I3_I0_int_0n[1], I26_c_0n[4], I26_I15_ha );
  OR2 I26_I15_I3_I0_I0 ( I26_c_0n[5], I26_I15_I3_I0_int_0n[0], I26_I15_I3_I0_int_0n[1] );
  AN2 I26_I16_I3_I0_I2 ( I26_I16_I3_I0_int_0n[0], I26_n_0n[5], I26_I16_I3_nsel_0n );
  AN2 I26_I16_I3_I0_I1 ( I26_I16_I3_I0_int_0n[1], I26_c_0n[5], I26_I16_ha );
  OR2 I26_I16_I3_I0_I0 ( I26_c_0n[6], I26_I16_I3_I0_int_0n[0], I26_I16_I3_I0_int_0n[1] );
  AN2 I26_I17_I3_I0_I2 ( I26_I17_I3_I0_int_0n[0], I26_n_0n[6], I26_I17_I3_nsel_0n );
  AN2 I26_I17_I3_I0_I1 ( I26_I17_I3_I0_int_0n[1], I26_c_0n[6], I26_I17_ha );
  OR2 I26_I17_I3_I0_I0 ( I26_c_0n[7], I26_I17_I3_I0_int_0n[0], I26_I17_I3_I0_int_0n[1] );
  AN2 I26_I18_I3_I0_I2 ( I26_I18_I3_I0_int_0n[0], I26_n_0n[7], I26_I18_I3_nsel_0n );
  AN2 I26_I18_I3_I0_I1 ( I26_I18_I3_I0_int_0n[1], I26_c_0n[7], I26_I18_ha );
  OR2 I26_I18_I3_I0_I0 ( I26_c_0n[8], I26_I18_I3_I0_int_0n[0], I26_I18_I3_I0_int_0n[1] );
endmodule

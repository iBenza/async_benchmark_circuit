
module Balsa_gcd16 ( activate_0r, activate_0a, x_0r, x_0a, x_0d, y_0r, y_0a, y_0d, z_0r, z_0a, z_0d, initialise );
  input [15:0] x_0d;
  input [15:0] y_0d;
  output [15:0] z_0d;
  input activate_0r, x_0a, y_0a, z_0a, initialise;
  output activate_0a, x_0r, y_0r, z_0r;

  wire activate_0r;
  wire activate_0a;
  wire x_0r;
  wire x_0a;
  wire [15:0] x_0d;
  wire y_0r;
  wire y_0a;
  wire [15:0] y_0d;
  wire z_0r;
  wire z_0a;
  wire [15:0] z_0d;
  wire initialise;
  wire c45_r;
  wire c45_a;
  wire [15:0] c45_d;
  wire c44_r;
  wire c44_a;
  wire [15:0] c44_d;
  wire c43_r;
  wire c42_r;
  wire c42_a;
  wire c40_a;
  wire c38_a;
  wire c37_r;
  wire c37_a;
  wire c36_r;
  wire c36_a;
  wire c36_d;
  wire [15:0] c34_d;
  wire c33_r;
  wire c33_d;
  wire c32_r;
  wire c32_d;
  wire c31_a;
  wire c30_a;
  wire c28_r;
  wire c27_r;
  wire [15:0] c24_d;
  wire c23_a;
  wire c22_r;
  wire c21_r;
  wire c20_r;
  wire c19_a;
  wire c18_a;
  wire [15:0] c18_d;
  wire [15:0] c15_d;
  wire c14_a;
  wire c13_r;
  wire c12_r;
  wire c11_r;
  wire c10_a;
  wire c9_a;
  wire [15:0] c9_d;
  wire I0_nbWriteReq_0n;
  wire I0_bWriteReq_0n;
  wire I0_nWriteReq_0n;
  wire I2_nbWriteReq_0n;
  wire I2_bWriteReq_0n;
  wire I2_nWriteReq_0n;
  wire I1_nselect_0n;
  wire I1_select_0n;
  wire I3_nselect_0n;
  wire I3_select_0n;
  wire I4_nReq_0n;
  wire I5_sreq_0n_1_;
  wire I5_I3_s;
  wire [1:0] I6_acks_0n;
  wire I6_I1_s_0n;
  wire I6_I2_s_0n;
  wire I9_nReq_0n;
  wire I9_guardAck_0n;
  wire I9_guardReq_0n;
  wire [15:0] I10_eq_0n;
  wire [3:0] I10_internal_0n;
  wire I9_I0_ns_0n;
  wire I11_I5_ns_0n;
  wire I15_nbWriteReq_0n;
  wire I15_bWriteReq_0n;
  wire I15_nWriteReq_0n;
  wire I16_vcc;
  wire I16_nxv_0n;
  wire I16_z_0n;
  wire I16_v_0n;
  wire [15:0] I16_n_0n;
  wire I16_addOut_0n_0_;
  wire I16_addOut_0n_1_;
  wire I16_addOut_0n_2_;
  wire I16_addOut_0n_3_;
  wire I16_addOut_0n_4_;
  wire I16_addOut_0n_5_;
  wire I16_addOut_0n_6_;
  wire I16_addOut_0n_7_;
  wire I16_addOut_0n_8_;
  wire I16_addOut_0n_9_;
  wire I16_addOut_0n_10_;
  wire I16_addOut_0n_11_;
  wire I16_addOut_0n_12_;
  wire I16_addOut_0n_13_;
  wire I16_addOut_0n_14_;
  wire I16_addOut_0n_15_;
  wire I16_c_0n_1_;
  wire I16_c_0n_2_;
  wire I16_c_0n_3_;
  wire I16_c_0n_4_;
  wire I16_c_0n_5_;
  wire I16_c_0n_6_;
  wire I16_c_0n_7_;
  wire I16_c_0n_8_;
  wire I16_c_0n_9_;
  wire I16_c_0n_10_;
  wire I16_c_0n_11_;
  wire I16_c_0n_12_;
  wire I16_c_0n_13_;
  wire I16_c_0n_14_;
  wire I16_c_0n_15_;
  wire I16_c_0n_16_;
  wire I16_nCv_0n_1_;
  wire I16_nCv_0n_2_;
  wire I16_nCv_0n_3_;
  wire I16_nCv_0n_4_;
  wire I16_nCv_0n_5_;
  wire I16_nCv_0n_6_;
  wire I16_nCv_0n_7_;
  wire I16_nCv_0n_8_;
  wire I16_nCv_0n_9_;
  wire I16_nCv_0n_10_;
  wire I16_nCv_0n_11_;
  wire I16_nCv_0n_12_;
  wire I16_nCv_0n_13_;
  wire I16_nCv_0n_14_;
  wire I16_nCv_0n_15_;
  wire I16_nCv_0n_16_;
  wire I16_nStart_0n;
  wire I16_start_0n;
  wire [7:0] I16_internal_0n;
  wire I5_I4_s_0n;
  wire I9_I1_s_0n;
  wire I12_I3_s_0n;
  wire I17_I3_s_0n;
  wire I22_I3_s_0n;
  wire I20_nbWriteReq_0n;
  wire I20_bWriteReq_0n;
  wire I20_nWriteReq_0n;
  wire I25_nbWriteReq_0n;
  wire I25_bWriteReq_0n;
  wire I25_nWriteReq_0n;
  wire I21_vcc;
  wire [15:0] I21_n_0n;
  wire [16:1] I21_c_0n;
  wire I21_nCv_0n_1_;
  wire I21_nCv_0n_2_;
  wire I21_nCv_0n_3_;
  wire I21_nCv_0n_4_;
  wire I21_nCv_0n_5_;
  wire I21_nCv_0n_6_;
  wire I21_nCv_0n_7_;
  wire I21_nCv_0n_8_;
  wire I21_nCv_0n_9_;
  wire I21_nCv_0n_10_;
  wire I21_nCv_0n_11_;
  wire I21_nCv_0n_12_;
  wire I21_nCv_0n_13_;
  wire I21_nCv_0n_14_;
  wire I21_nCv_0n_15_;
  wire I21_nCv_0n_16_;
  wire I21_nStart_0n;
  wire I21_start_0n;
  wire [3:0] I21_internal_0n;
  wire I26_vcc;
  wire [15:0] I26_n_0n;
  wire [16:1] I26_c_0n;
  wire I26_nCv_0n_1_;
  wire I26_nCv_0n_2_;
  wire I26_nCv_0n_3_;
  wire I26_nCv_0n_4_;
  wire I26_nCv_0n_5_;
  wire I26_nCv_0n_6_;
  wire I26_nCv_0n_7_;
  wire I26_nCv_0n_8_;
  wire I26_nCv_0n_9_;
  wire I26_nCv_0n_10_;
  wire I26_nCv_0n_11_;
  wire I26_nCv_0n_12_;
  wire I26_nCv_0n_13_;
  wire I26_nCv_0n_14_;
  wire I26_nCv_0n_15_;
  wire I26_nCv_0n_16_;
  wire I26_nStart_0n;
  wire I26_start_0n;
  wire [3:0] I26_internal_0n;
  wire I16_I13_cv;
  wire I16_I13_ha;
  wire I16_I13_start;
  wire I16_I14_cv;
  wire I16_I14_ha;
  wire I16_I14_start;
  wire I16_I15_cv;
  wire I16_I15_ha;
  wire I16_I15_start;
  wire I16_I16_cv;
  wire I16_I16_ha;
  wire I16_I16_start;
  wire I16_I17_cv;
  wire I16_I17_ha;
  wire I16_I17_start;
  wire I16_I18_cv;
  wire I16_I18_ha;
  wire I16_I18_start;
  wire I16_I19_cv;
  wire I16_I19_ha;
  wire I16_I19_start;
  wire I16_I20_cv;
  wire I16_I20_ha;
  wire I16_I20_start;
  wire I16_I21_cv;
  wire I16_I21_ha;
  wire I16_I21_start;
  wire I16_I22_cv;
  wire I16_I22_ha;
  wire I16_I22_start;
  wire I16_I23_cv;
  wire I16_I23_ha;
  wire I16_I23_start;
  wire I16_I24_cv;
  wire I16_I24_ha;
  wire I16_I24_start;
  wire I16_I25_cv;
  wire I16_I25_ha;
  wire I16_I25_start;
  wire I16_I26_cv;
  wire I16_I26_ha;
  wire I16_I26_start;
  wire I16_I27_cv;
  wire I16_I27_ha;
  wire I16_I27_start;
  wire I16_I28_cv;
  wire I16_I28_ha;
  wire I16_I28_start;
  wire I21_I21_cv;
  wire I21_I21_ha;
  wire I21_I21_start;
  wire I21_I22_cv;
  wire I21_I22_ha;
  wire I21_I22_start;
  wire I21_I23_cv;
  wire I21_I23_ha;
  wire I21_I23_start;
  wire I21_I24_cv;
  wire I21_I24_ha;
  wire I21_I24_start;
  wire I21_I25_cv;
  wire I21_I25_ha;
  wire I21_I25_start;
  wire I21_I26_cv;
  wire I21_I26_ha;
  wire I21_I26_start;
  wire I21_I27_cv;
  wire I21_I27_ha;
  wire I21_I27_start;
  wire I21_I28_cv;
  wire I21_I28_ha;
  wire I21_I28_start;
  wire I21_I29_cv;
  wire I21_I29_ha;
  wire I21_I29_start;
  wire I21_I30_cv;
  wire I21_I30_ha;
  wire I21_I30_start;
  wire I21_I31_cv;
  wire I21_I31_ha;
  wire I21_I31_start;
  wire I21_I32_cv;
  wire I21_I32_ha;
  wire I21_I32_start;
  wire I21_I33_cv;
  wire I21_I33_ha;
  wire I21_I33_start;
  wire I21_I34_cv;
  wire I21_I34_ha;
  wire I21_I34_start;
  wire I21_I35_cv;
  wire I21_I35_ha;
  wire I21_I35_start;
  wire I21_I36_cv;
  wire I21_I36_ha;
  wire I21_I36_start;
  wire I26_I21_cv;
  wire I26_I21_ha;
  wire I26_I21_start;
  wire I26_I22_cv;
  wire I26_I22_ha;
  wire I26_I22_start;
  wire I26_I23_cv;
  wire I26_I23_ha;
  wire I26_I23_start;
  wire I26_I24_cv;
  wire I26_I24_ha;
  wire I26_I24_start;
  wire I26_I25_cv;
  wire I26_I25_ha;
  wire I26_I25_start;
  wire I26_I26_cv;
  wire I26_I26_ha;
  wire I26_I26_start;
  wire I26_I27_cv;
  wire I26_I27_ha;
  wire I26_I27_start;
  wire I26_I28_cv;
  wire I26_I28_ha;
  wire I26_I28_start;
  wire I26_I29_cv;
  wire I26_I29_ha;
  wire I26_I29_start;
  wire I26_I30_cv;
  wire I26_I30_ha;
  wire I26_I30_start;
  wire I26_I31_cv;
  wire I26_I31_ha;
  wire I26_I31_start;
  wire I26_I32_cv;
  wire I26_I32_ha;
  wire I26_I32_start;
  wire I26_I33_cv;
  wire I26_I33_ha;
  wire I26_I33_start;
  wire I26_I34_cv;
  wire I26_I34_ha;
  wire I26_I34_start;
  wire I26_I35_cv;
  wire I26_I35_ha;
  wire I26_I35_start;
  wire I26_I36_cv;
  wire I26_I36_ha;
  wire I26_I36_start;
  wire I16_I13_I2_nsel_0n;
  wire I16_I14_I2_nsel_0n;
  wire I16_I15_I2_nsel_0n;
  wire I16_I16_I2_nsel_0n;
  wire I16_I17_I2_nsel_0n;
  wire I16_I18_I2_nsel_0n;
  wire I16_I19_I2_nsel_0n;
  wire I16_I20_I2_nsel_0n;
  wire I16_I21_I2_nsel_0n;
  wire I16_I22_I2_nsel_0n;
  wire I16_I23_I2_nsel_0n;
  wire I16_I24_I2_nsel_0n;
  wire I16_I25_I2_nsel_0n;
  wire I16_I26_I2_nsel_0n;
  wire I16_I27_I2_nsel_0n;
  wire I16_I28_I2_nsel_0n;
  wire I21_I21_I2_nsel_0n;
  wire I21_I22_I2_nsel_0n;
  wire I21_I23_I2_nsel_0n;
  wire I21_I24_I2_nsel_0n;
  wire I21_I25_I2_nsel_0n;
  wire I21_I26_I2_nsel_0n;
  wire I21_I27_I2_nsel_0n;
  wire I21_I28_I2_nsel_0n;
  wire I21_I29_I2_nsel_0n;
  wire I21_I30_I2_nsel_0n;
  wire I21_I31_I2_nsel_0n;
  wire I21_I32_I2_nsel_0n;
  wire I21_I33_I2_nsel_0n;
  wire I21_I34_I2_nsel_0n;
  wire I21_I35_I2_nsel_0n;
  wire I21_I36_I2_nsel_0n;
  wire I26_I21_I2_nsel_0n;
  wire I26_I22_I2_nsel_0n;
  wire I26_I23_I2_nsel_0n;
  wire I26_I24_I2_nsel_0n;
  wire I26_I25_I2_nsel_0n;
  wire I26_I26_I2_nsel_0n;
  wire I26_I27_I2_nsel_0n;
  wire I26_I28_I2_nsel_0n;
  wire I26_I29_I2_nsel_0n;
  wire I26_I30_I2_nsel_0n;
  wire I26_I31_I2_nsel_0n;
  wire I26_I32_I2_nsel_0n;
  wire I26_I33_I2_nsel_0n;
  wire I26_I34_I2_nsel_0n;
  wire I26_I35_I2_nsel_0n;
  wire I26_I36_I2_nsel_0n;
  wire [1:0] I16_I13_I2_I0_int_0n;
  wire [1:0] I16_I14_I2_I0_int_0n;
  wire [1:0] I16_I15_I2_I0_int_0n;
  wire [1:0] I16_I16_I2_I0_int_0n;
  wire [1:0] I16_I17_I2_I0_int_0n;
  wire [1:0] I16_I18_I2_I0_int_0n;
  wire [1:0] I16_I19_I2_I0_int_0n;
  wire [1:0] I16_I20_I2_I0_int_0n;
  wire [1:0] I16_I21_I2_I0_int_0n;
  wire [1:0] I16_I22_I2_I0_int_0n;
  wire [1:0] I16_I23_I2_I0_int_0n;
  wire [1:0] I16_I24_I2_I0_int_0n;
  wire [1:0] I16_I25_I2_I0_int_0n;
  wire [1:0] I16_I26_I2_I0_int_0n;
  wire [1:0] I16_I27_I2_I0_int_0n;
  wire [1:0] I16_I28_I2_I0_int_0n;
  wire [1:0] I21_I21_I2_I0_int_0n;
  wire [1:0] I21_I22_I2_I0_int_0n;
  wire [1:0] I21_I23_I2_I0_int_0n;
  wire [1:0] I21_I24_I2_I0_int_0n;
  wire [1:0] I21_I25_I2_I0_int_0n;
  wire [1:0] I21_I26_I2_I0_int_0n;
  wire [1:0] I21_I27_I2_I0_int_0n;
  wire [1:0] I21_I28_I2_I0_int_0n;
  wire [1:0] I21_I29_I2_I0_int_0n;
  wire [1:0] I21_I30_I2_I0_int_0n;
  wire [1:0] I21_I31_I2_I0_int_0n;
  wire [1:0] I21_I32_I2_I0_int_0n;
  wire [1:0] I21_I33_I2_I0_int_0n;
  wire [1:0] I21_I34_I2_I0_int_0n;
  wire [1:0] I21_I35_I2_I0_int_0n;
  wire [1:0] I21_I36_I2_I0_int_0n;
  wire [1:0] I26_I21_I2_I0_int_0n;
  wire [1:0] I26_I22_I2_I0_int_0n;
  wire [1:0] I26_I23_I2_I0_int_0n;
  wire [1:0] I26_I24_I2_I0_int_0n;
  wire [1:0] I26_I25_I2_I0_int_0n;
  wire [1:0] I26_I26_I2_I0_int_0n;
  wire [1:0] I26_I27_I2_I0_int_0n;
  wire [1:0] I26_I28_I2_I0_int_0n;
  wire [1:0] I26_I29_I2_I0_int_0n;
  wire [1:0] I26_I30_I2_I0_int_0n;
  wire [1:0] I26_I31_I2_I0_int_0n;
  wire [1:0] I26_I32_I2_I0_int_0n;
  wire [1:0] I26_I33_I2_I0_int_0n;
  wire [1:0] I26_I34_I2_I0_int_0n;
  wire [1:0] I26_I35_I2_I0_int_0n;
  wire [1:0] I26_I36_I2_I0_int_0n;
  wire I1_I0_nsel_0n;
  wire I1_I1_nsel_0n;
  wire I1_I2_nsel_0n;
  wire I1_I3_nsel_0n;
  wire I1_I4_nsel_0n;
  wire I1_I5_nsel_0n;
  wire I1_I6_nsel_0n;
  wire I1_I7_nsel_0n;
  wire I1_I8_nsel_0n;
  wire I1_I9_nsel_0n;
  wire I1_I10_nsel_0n;
  wire I1_I11_nsel_0n;
  wire I1_I12_nsel_0n;
  wire I1_I13_nsel_0n;
  wire I1_I14_nsel_0n;
  wire I1_I15_nsel_0n;
  wire I1_I16_nsel_0n;
  wire I3_I0_nsel_0n;
  wire I3_I1_nsel_0n;
  wire I3_I2_nsel_0n;
  wire I3_I3_nsel_0n;
  wire I3_I4_nsel_0n;
  wire I3_I5_nsel_0n;
  wire I3_I6_nsel_0n;
  wire I3_I7_nsel_0n;
  wire I3_I8_nsel_0n;
  wire I3_I9_nsel_0n;
  wire I3_I10_nsel_0n;
  wire I3_I11_nsel_0n;
  wire I3_I12_nsel_0n;
  wire I3_I13_nsel_0n;
  wire I3_I14_nsel_0n;
  wire I3_I15_nsel_0n;
  wire I3_I16_nsel_0n;
  wire I16_I13_I3_nsel_0n;
  wire I16_I14_I3_nsel_0n;
  wire I16_I15_I3_nsel_0n;
  wire I16_I16_I3_nsel_0n;
  wire I16_I17_I3_nsel_0n;
  wire I16_I18_I3_nsel_0n;
  wire I16_I19_I3_nsel_0n;
  wire I16_I20_I3_nsel_0n;
  wire I16_I21_I3_nsel_0n;
  wire I16_I22_I3_nsel_0n;
  wire I16_I23_I3_nsel_0n;
  wire I16_I24_I3_nsel_0n;
  wire I16_I25_I3_nsel_0n;
  wire I16_I26_I3_nsel_0n;
  wire I16_I27_I3_nsel_0n;
  wire I16_I28_I3_nsel_0n;
  wire I21_I21_I3_nsel_0n;
  wire I21_I22_I3_nsel_0n;
  wire I21_I23_I3_nsel_0n;
  wire I21_I24_I3_nsel_0n;
  wire I21_I25_I3_nsel_0n;
  wire I21_I26_I3_nsel_0n;
  wire I21_I27_I3_nsel_0n;
  wire I21_I28_I3_nsel_0n;
  wire I21_I29_I3_nsel_0n;
  wire I21_I30_I3_nsel_0n;
  wire I21_I31_I3_nsel_0n;
  wire I21_I32_I3_nsel_0n;
  wire I21_I33_I3_nsel_0n;
  wire I21_I34_I3_nsel_0n;
  wire I21_I35_I3_nsel_0n;
  wire I21_I36_I3_nsel_0n;
  wire I26_I21_I3_nsel_0n;
  wire I26_I22_I3_nsel_0n;
  wire I26_I23_I3_nsel_0n;
  wire I26_I24_I3_nsel_0n;
  wire I26_I25_I3_nsel_0n;
  wire I26_I26_I3_nsel_0n;
  wire I26_I27_I3_nsel_0n;
  wire I26_I28_I3_nsel_0n;
  wire I26_I29_I3_nsel_0n;
  wire I26_I30_I3_nsel_0n;
  wire I26_I31_I3_nsel_0n;
  wire I26_I32_I3_nsel_0n;
  wire I26_I33_I3_nsel_0n;
  wire I26_I34_I3_nsel_0n;
  wire I26_I35_I3_nsel_0n;
  wire I26_I36_I3_nsel_0n;
  wire [1:0] I1_I0_I0_int_0n;
  wire [1:0] I1_I1_I0_int_0n;
  wire [1:0] I1_I2_I0_int_0n;
  wire [1:0] I1_I3_I0_int_0n;
  wire [1:0] I1_I4_I0_int_0n;
  wire [1:0] I1_I5_I0_int_0n;
  wire [1:0] I1_I6_I0_int_0n;
  wire [1:0] I1_I7_I0_int_0n;
  wire [1:0] I1_I8_I0_int_0n;
  wire [1:0] I1_I9_I0_int_0n;
  wire [1:0] I1_I10_I0_int_0n;
  wire [1:0] I1_I11_I0_int_0n;
  wire [1:0] I1_I12_I0_int_0n;
  wire [1:0] I1_I13_I0_int_0n;
  wire [1:0] I1_I14_I0_int_0n;
  wire [1:0] I1_I15_I0_int_0n;
  wire [1:0] I1_I16_I0_int_0n;
  wire [1:0] I3_I0_I0_int_0n;
  wire [1:0] I3_I1_I0_int_0n;
  wire [1:0] I3_I2_I0_int_0n;
  wire [1:0] I3_I3_I0_int_0n;
  wire [1:0] I3_I4_I0_int_0n;
  wire [1:0] I3_I5_I0_int_0n;
  wire [1:0] I3_I6_I0_int_0n;
  wire [1:0] I3_I7_I0_int_0n;
  wire [1:0] I3_I8_I0_int_0n;
  wire [1:0] I3_I9_I0_int_0n;
  wire [1:0] I3_I10_I0_int_0n;
  wire [1:0] I3_I11_I0_int_0n;
  wire [1:0] I3_I12_I0_int_0n;
  wire [1:0] I3_I13_I0_int_0n;
  wire [1:0] I3_I14_I0_int_0n;
  wire [1:0] I3_I15_I0_int_0n;
  wire [1:0] I3_I16_I0_int_0n;
  wire [1:0] I16_I13_I3_I0_int_0n;
  wire [1:0] I16_I14_I3_I0_int_0n;
  wire [1:0] I16_I15_I3_I0_int_0n;
  wire [1:0] I16_I16_I3_I0_int_0n;
  wire [1:0] I16_I17_I3_I0_int_0n;
  wire [1:0] I16_I18_I3_I0_int_0n;
  wire [1:0] I16_I19_I3_I0_int_0n;
  wire [1:0] I16_I20_I3_I0_int_0n;
  wire [1:0] I16_I21_I3_I0_int_0n;
  wire [1:0] I16_I22_I3_I0_int_0n;
  wire [1:0] I16_I23_I3_I0_int_0n;
  wire [1:0] I16_I24_I3_I0_int_0n;
  wire [1:0] I16_I25_I3_I0_int_0n;
  wire [1:0] I16_I26_I3_I0_int_0n;
  wire [1:0] I16_I27_I3_I0_int_0n;
  wire [1:0] I16_I28_I3_I0_int_0n;
  wire [1:0] I21_I21_I3_I0_int_0n;
  wire [1:0] I21_I22_I3_I0_int_0n;
  wire [1:0] I21_I23_I3_I0_int_0n;
  wire [1:0] I21_I24_I3_I0_int_0n;
  wire [1:0] I21_I25_I3_I0_int_0n;
  wire [1:0] I21_I26_I3_I0_int_0n;
  wire [1:0] I21_I27_I3_I0_int_0n;
  wire [1:0] I21_I28_I3_I0_int_0n;
  wire [1:0] I21_I29_I3_I0_int_0n;
  wire [1:0] I21_I30_I3_I0_int_0n;
  wire [1:0] I21_I31_I3_I0_int_0n;
  wire [1:0] I21_I32_I3_I0_int_0n;
  wire [1:0] I21_I33_I3_I0_int_0n;
  wire [1:0] I21_I34_I3_I0_int_0n;
  wire [1:0] I21_I35_I3_I0_int_0n;
  wire [1:0] I21_I36_I3_I0_int_0n;
  wire [1:0] I26_I21_I3_I0_int_0n;
  wire [1:0] I26_I22_I3_I0_int_0n;
  wire [1:0] I26_I23_I3_I0_int_0n;
  wire [1:0] I26_I24_I3_I0_int_0n;
  wire [1:0] I26_I25_I3_I0_int_0n;
  wire [1:0] I26_I26_I3_I0_int_0n;
  wire [1:0] I26_I27_I3_I0_int_0n;
  wire [1:0] I26_I28_I3_I0_int_0n;
  wire [1:0] I26_I29_I3_I0_int_0n;
  wire [1:0] I26_I30_I3_I0_int_0n;
  wire [1:0] I26_I31_I3_I0_int_0n;
  wire [1:0] I26_I32_I3_I0_int_0n;
  wire [1:0] I26_I33_I3_I0_int_0n;
  wire [1:0] I26_I34_I3_I0_int_0n;
  wire [1:0] I26_I35_I3_I0_int_0n;
  wire [1:0] I26_I36_I3_I0_int_0n;

  IV I0_I104 ( I0_nWriteReq_0n, c45_r );
  IV I0_I103 ( I0_bWriteReq_0n, I0_nWriteReq_0n );
  IV I0_I102 ( I0_nbWriteReq_0n, I0_bWriteReq_0n );
  IV I0_I101 ( c45_a, I0_nbWriteReq_0n );
  LD1 I0_I100 ( c45_d[15], I0_bWriteReq_0n, z_0d[15] );
  LD1 I0_I99 ( c45_d[14], I0_bWriteReq_0n, z_0d[14] );
  LD1 I0_I98 ( c45_d[13], I0_bWriteReq_0n, z_0d[13] );
  LD1 I0_I97 ( c45_d[12], I0_bWriteReq_0n, z_0d[12] );
  LD1 I0_I96 ( c45_d[11], I0_bWriteReq_0n, z_0d[11] );
  LD1 I0_I95 ( c45_d[10], I0_bWriteReq_0n, z_0d[10] );
  LD1 I0_I94 ( c45_d[9], I0_bWriteReq_0n, z_0d[9] );
  LD1 I0_I93 ( c45_d[8], I0_bWriteReq_0n, z_0d[8] );
  LD1 I0_I92 ( c45_d[7], I0_bWriteReq_0n, z_0d[7] );
  LD1 I0_I91 ( c45_d[6], I0_bWriteReq_0n, z_0d[6] );
  LD1 I0_I90 ( c45_d[5], I0_bWriteReq_0n, z_0d[5] );
  LD1 I0_I89 ( c45_d[4], I0_bWriteReq_0n, z_0d[4] );
  LD1 I0_I88 ( c45_d[3], I0_bWriteReq_0n, z_0d[3] );
  LD1 I0_I87 ( c45_d[2], I0_bWriteReq_0n, z_0d[2] );
  LD1 I0_I86 ( c45_d[1], I0_bWriteReq_0n, z_0d[1] );
  LD1 I0_I85 ( c45_d[0], I0_bWriteReq_0n, z_0d[0] );
  IV I2_I87 ( I2_nWriteReq_0n, c44_r );
  IV I2_I86 ( I2_bWriteReq_0n, I2_nWriteReq_0n );
  IV I2_I85 ( I2_nbWriteReq_0n, I2_bWriteReq_0n );
  IV I2_I84 ( c44_a, I2_nbWriteReq_0n );
  LD1 I2_I83 ( c44_d[15], I2_bWriteReq_0n, c34_d[15] );
  LD1 I2_I82 ( c44_d[14], I2_bWriteReq_0n, c34_d[14] );
  LD1 I2_I81 ( c44_d[13], I2_bWriteReq_0n, c34_d[13] );
  LD1 I2_I80 ( c44_d[12], I2_bWriteReq_0n, c34_d[12] );
  LD1 I2_I79 ( c44_d[11], I2_bWriteReq_0n, c34_d[11] );
  LD1 I2_I78 ( c44_d[10], I2_bWriteReq_0n, c34_d[10] );
  LD1 I2_I77 ( c44_d[9], I2_bWriteReq_0n, c34_d[9] );
  LD1 I2_I76 ( c44_d[8], I2_bWriteReq_0n, c34_d[8] );
  LD1 I2_I75 ( c44_d[7], I2_bWriteReq_0n, c34_d[7] );
  LD1 I2_I74 ( c44_d[6], I2_bWriteReq_0n, c34_d[6] );
  LD1 I2_I73 ( c44_d[5], I2_bWriteReq_0n, c34_d[5] );
  LD1 I2_I72 ( c44_d[4], I2_bWriteReq_0n, c34_d[4] );
  LD1 I2_I71 ( c44_d[3], I2_bWriteReq_0n, c34_d[3] );
  LD1 I2_I70 ( c44_d[2], I2_bWriteReq_0n, c34_d[2] );
  LD1 I2_I69 ( c44_d[1], I2_bWriteReq_0n, c34_d[1] );
  LD1 I2_I68 ( c44_d[0], I2_bWriteReq_0n, c34_d[0] );
  SRFF I1_I19 ( x_0a, c22_r, I1_select_0n, I1_nselect_0n );
  AN2 I1_I18 ( c40_a, I1_select_0n, c45_a );
  AN2 I1_I17 ( c19_a, I1_nselect_0n, c45_a );
  SRFF I3_I19 ( y_0a, c13_r, I3_select_0n, I3_nselect_0n );
  AN2 I3_I18 ( c38_a, I3_select_0n, c44_a );
  AN2 I3_I17 ( c10_a, I3_nselect_0n, c44_a );
  NR2 I4_I1 ( c43_r, I4_nReq_0n, z_0a );
  IV I4_I0 ( I4_nReq_0n, activate_0r );
  GND I4_gnd_cell_instance ( activate_0a );
  C2R I5_I3_I2 ( z_0r, c37_a, I5_sreq_0n_1_, initialise );
  IV I5_I3_I1 ( I5_I3_s, z_0r );
  AN2 I5_I3_I0 ( c37_r, I5_sreq_0n_1_, I5_I3_s );
  C2 I6_I0 ( c42_a, I6_acks_0n[0], I6_acks_0n[1] );
  AN2 I6_I1_I2 ( x_0r, c42_r, I6_I1_s_0n );
  IV I6_I1_I1 ( I6_I1_s_0n, I6_acks_0n[0] );
  ACU0D1 I6_I1_I0 ( I6_acks_0n[0], c40_a, c42_r );
  AN2 I6_I2_I2 ( y_0r, c42_r, I6_I2_s_0n );
  IV I6_I2_I1 ( I6_I2_s_0n, I6_acks_0n[1] );
  ACU0D1 I6_I2_I0 ( I6_acks_0n[1], c38_a, c42_r );
  NR2 I9_I3 ( I9_guardReq_0n, I9_nReq_0n, c31_a );
  IV I9_I2 ( I9_nReq_0n, c37_r );
  C2 I10_I55 ( c36_a, c36_r, c36_r );
  EO I10_I20 ( I10_eq_0n[15], z_0d[15], c34_d[15] );
  EO I10_I19 ( I10_eq_0n[14], z_0d[14], c34_d[14] );
  EO I10_I18 ( I10_eq_0n[13], z_0d[13], c34_d[13] );
  EO I10_I17 ( I10_eq_0n[12], z_0d[12], c34_d[12] );
  EO I10_I16 ( I10_eq_0n[11], z_0d[11], c34_d[11] );
  EO I10_I15 ( I10_eq_0n[10], z_0d[10], c34_d[10] );
  EO I10_I14 ( I10_eq_0n[9], z_0d[9], c34_d[9] );
  EO I10_I13 ( I10_eq_0n[8], z_0d[8], c34_d[8] );
  EO I10_I12 ( I10_eq_0n[7], z_0d[7], c34_d[7] );
  EO I10_I11 ( I10_eq_0n[6], z_0d[6], c34_d[6] );
  EO I10_I10 ( I10_eq_0n[5], z_0d[5], c34_d[5] );
  EO I10_I9 ( I10_eq_0n[4], z_0d[4], c34_d[4] );
  EO I10_I8 ( I10_eq_0n[3], z_0d[3], c34_d[3] );
  EO I10_I7 ( I10_eq_0n[2], z_0d[2], c34_d[2] );
  EO I10_I6 ( I10_eq_0n[1], z_0d[1], c34_d[1] );
  EO I10_I5 ( I10_eq_0n[0], z_0d[0], c34_d[0] );
  ND4 I10_I4 ( c36_d, I10_internal_0n[0], I10_internal_0n[1], I10_internal_0n[2], I10_internal_0n[3] );
  NR4 I10_I3 ( I10_internal_0n[3], I10_eq_0n[12], I10_eq_0n[13], I10_eq_0n[14], I10_eq_0n[15] );
  NR4 I10_I2 ( I10_internal_0n[2], I10_eq_0n[8], I10_eq_0n[9], I10_eq_0n[10], I10_eq_0n[11] );
  NR4 I10_I1 ( I10_internal_0n[1], I10_eq_0n[4], I10_eq_0n[5], I10_eq_0n[6], I10_eq_0n[7] );
  NR4 I10_I0 ( I10_internal_0n[0], I10_eq_0n[0], I10_eq_0n[1], I10_eq_0n[2], I10_eq_0n[3] );
  OR2 I11_I0 ( c31_a, c10_a, c19_a );
  IV I9_I0_I2 ( I9_I0_ns_0n, c36_d );
  AN2 I9_I0_I1 ( c37_a, c36_a, I9_I0_ns_0n );
  AN2 I9_I0_I0 ( I9_guardAck_0n, c36_a, c36_d );
  IV I11_I5_I2 ( I11_I5_ns_0n, c33_d );
  AN2 I11_I5_I1 ( c11_r, c33_r, I11_I5_ns_0n );
  AN2 I11_I5_I0 ( c20_r, c33_r, c33_d );
  IV I15_I6 ( I15_nWriteReq_0n, c32_r );
  IV I15_I5 ( I15_bWriteReq_0n, I15_nWriteReq_0n );
  IV I15_I4 ( I15_nbWriteReq_0n, I15_bWriteReq_0n );
  IV I15_I3 ( c30_a, I15_nbWriteReq_0n );
  LD1 I15_I2 ( c32_d, I15_bWriteReq_0n, c33_d );
  C2 I16_I65 ( I16_start_0n, c27_r, c27_r );
  IV I16_I47 ( I16_n_0n[15], c34_d[15] );
  IV I16_I46 ( I16_n_0n[14], c34_d[14] );
  IV I16_I45 ( I16_n_0n[13], c34_d[13] );
  IV I16_I44 ( I16_n_0n[12], c34_d[12] );
  IV I16_I43 ( I16_n_0n[11], c34_d[11] );
  IV I16_I42 ( I16_n_0n[10], c34_d[10] );
  IV I16_I41 ( I16_n_0n[9], c34_d[9] );
  IV I16_I40 ( I16_n_0n[8], c34_d[8] );
  IV I16_I39 ( I16_n_0n[7], c34_d[7] );
  IV I16_I38 ( I16_n_0n[6], c34_d[6] );
  IV I16_I37 ( I16_n_0n[5], c34_d[5] );
  IV I16_I36 ( I16_n_0n[4], c34_d[4] );
  IV I16_I35 ( I16_n_0n[3], c34_d[3] );
  IV I16_I34 ( I16_n_0n[2], c34_d[2] );
  IV I16_I33 ( I16_n_0n[1], c34_d[1] );
  IV I16_I32 ( I16_n_0n[0], c34_d[0] );
  IV I16_I31 ( I16_nStart_0n, I16_start_0n );
  EO I16_I12 ( I16_v_0n, I16_c_0n_15_, I16_c_0n_16_ );
  AN4 I16_I11 ( c32_r, I16_internal_0n[4], I16_internal_0n[5], I16_internal_0n[6], I16_internal_0n[7] );
  NR4 I16_I10 ( I16_internal_0n[7], I16_nCv_0n_13_, I16_nCv_0n_14_, I16_nCv_0n_15_, I16_nCv_0n_16_ );
  NR4 I16_I9 ( I16_internal_0n[6], I16_nCv_0n_9_, I16_nCv_0n_10_, I16_nCv_0n_11_, I16_nCv_0n_12_ );
  NR4 I16_I8 ( I16_internal_0n[5], I16_nCv_0n_5_, I16_nCv_0n_6_, I16_nCv_0n_7_, I16_nCv_0n_8_ );
  NR4 I16_I7 ( I16_internal_0n[4], I16_nCv_0n_1_, I16_nCv_0n_2_, I16_nCv_0n_3_, I16_nCv_0n_4_ );
  AN4 I16_I6 ( I16_z_0n, I16_internal_0n[0], I16_internal_0n[1], I16_internal_0n[2], I16_internal_0n[3] );
  NR4 I16_I5 ( I16_internal_0n[3], I16_addOut_0n_12_, I16_addOut_0n_13_, I16_addOut_0n_14_, I16_addOut_0n_15_ );
  NR4 I16_I4 ( I16_internal_0n[2], I16_addOut_0n_8_, I16_addOut_0n_9_, I16_addOut_0n_10_, I16_addOut_0n_11_ );
  NR4 I16_I3 ( I16_internal_0n[1], I16_addOut_0n_4_, I16_addOut_0n_5_, I16_addOut_0n_6_, I16_addOut_0n_7_ );
  NR4 I16_I2 ( I16_internal_0n[0], I16_addOut_0n_0_, I16_addOut_0n_1_, I16_addOut_0n_2_, I16_addOut_0n_3_ );
  EO I16_I1 ( I16_nxv_0n, I16_v_0n, I16_addOut_0n_15_ );
  NR2 I16_I0 ( c32_d, I16_z_0n, I16_nxv_0n );
  VCC I16_vcc_cell_instance ( I16_vcc );
  AN2 I5_I4_I2 ( c42_r, c43_r, I5_I4_s_0n );
  NR2 I5_I4_I1 ( I5_sreq_0n_1_, c42_a, I5_I4_s_0n );
  NC2P I5_I4_I0 ( I5_I4_s_0n, c43_r, c42_a );
  AN2 I9_I1_I2 ( c36_r, I9_guardReq_0n, I9_I1_s_0n );
  NR2 I9_I1_I1 ( c28_r, I9_guardAck_0n, I9_I1_s_0n );
  NC2P I9_I1_I0 ( I9_I1_s_0n, I9_guardReq_0n, I9_guardAck_0n );
  AN2 I12_I3_I2 ( c27_r, c28_r, I12_I3_s_0n );
  NR2 I12_I3_I1 ( c33_r, c30_a, I12_I3_s_0n );
  NC2P I12_I3_I0 ( I12_I3_s_0n, c28_r, c30_a );
  AN2 I17_I3_I2 ( c21_r, c20_r, I17_I3_s_0n );
  NR2 I17_I3_I1 ( c22_r, c23_a, I17_I3_s_0n );
  NC2P I17_I3_I0 ( I17_I3_s_0n, c20_r, c23_a );
  AN2 I22_I3_I2 ( c12_r, c11_r, I22_I3_s_0n );
  NR2 I22_I3_I1 ( c13_r, c14_a, I22_I3_s_0n );
  NC2P I22_I3_I0 ( I22_I3_s_0n, c11_r, c14_a );
  IV I20_I36 ( I20_nWriteReq_0n, c18_a );
  IV I20_I35 ( I20_bWriteReq_0n, I20_nWriteReq_0n );
  IV I20_I34 ( I20_nbWriteReq_0n, I20_bWriteReq_0n );
  IV I20_I33 ( c23_a, I20_nbWriteReq_0n );
  LD1 I20_I32 ( c18_d[15], I20_bWriteReq_0n, c24_d[15] );
  LD1 I20_I31 ( c18_d[14], I20_bWriteReq_0n, c24_d[14] );
  LD1 I20_I30 ( c18_d[13], I20_bWriteReq_0n, c24_d[13] );
  LD1 I20_I29 ( c18_d[12], I20_bWriteReq_0n, c24_d[12] );
  LD1 I20_I28 ( c18_d[11], I20_bWriteReq_0n, c24_d[11] );
  LD1 I20_I27 ( c18_d[10], I20_bWriteReq_0n, c24_d[10] );
  LD1 I20_I26 ( c18_d[9], I20_bWriteReq_0n, c24_d[9] );
  LD1 I20_I25 ( c18_d[8], I20_bWriteReq_0n, c24_d[8] );
  LD1 I20_I24 ( c18_d[7], I20_bWriteReq_0n, c24_d[7] );
  LD1 I20_I23 ( c18_d[6], I20_bWriteReq_0n, c24_d[6] );
  LD1 I20_I22 ( c18_d[5], I20_bWriteReq_0n, c24_d[5] );
  LD1 I20_I21 ( c18_d[4], I20_bWriteReq_0n, c24_d[4] );
  LD1 I20_I20 ( c18_d[3], I20_bWriteReq_0n, c24_d[3] );
  LD1 I20_I19 ( c18_d[2], I20_bWriteReq_0n, c24_d[2] );
  LD1 I20_I18 ( c18_d[1], I20_bWriteReq_0n, c24_d[1] );
  LD1 I20_I17 ( c18_d[0], I20_bWriteReq_0n, c24_d[0] );
  IV I25_I36 ( I25_nWriteReq_0n, c9_a );
  IV I25_I35 ( I25_bWriteReq_0n, I25_nWriteReq_0n );
  IV I25_I34 ( I25_nbWriteReq_0n, I25_bWriteReq_0n );
  IV I25_I33 ( c14_a, I25_nbWriteReq_0n );
  LD1 I25_I32 ( c9_d[15], I25_bWriteReq_0n, c15_d[15] );
  LD1 I25_I31 ( c9_d[14], I25_bWriteReq_0n, c15_d[14] );
  LD1 I25_I30 ( c9_d[13], I25_bWriteReq_0n, c15_d[13] );
  LD1 I25_I29 ( c9_d[12], I25_bWriteReq_0n, c15_d[12] );
  LD1 I25_I28 ( c9_d[11], I25_bWriteReq_0n, c15_d[11] );
  LD1 I25_I27 ( c9_d[10], I25_bWriteReq_0n, c15_d[10] );
  LD1 I25_I26 ( c9_d[9], I25_bWriteReq_0n, c15_d[9] );
  LD1 I25_I25 ( c9_d[8], I25_bWriteReq_0n, c15_d[8] );
  LD1 I25_I24 ( c9_d[7], I25_bWriteReq_0n, c15_d[7] );
  LD1 I25_I23 ( c9_d[6], I25_bWriteReq_0n, c15_d[6] );
  LD1 I25_I22 ( c9_d[5], I25_bWriteReq_0n, c15_d[5] );
  LD1 I25_I21 ( c9_d[4], I25_bWriteReq_0n, c15_d[4] );
  LD1 I25_I20 ( c9_d[3], I25_bWriteReq_0n, c15_d[3] );
  LD1 I25_I19 ( c9_d[2], I25_bWriteReq_0n, c15_d[2] );
  LD1 I25_I18 ( c9_d[1], I25_bWriteReq_0n, c15_d[1] );
  LD1 I25_I17 ( c9_d[0], I25_bWriteReq_0n, c15_d[0] );
  C2 I21_I73 ( I21_start_0n, c21_r, c21_r );
  IV I21_I55 ( I21_n_0n[15], c34_d[15] );
  IV I21_I54 ( I21_n_0n[14], c34_d[14] );
  IV I21_I53 ( I21_n_0n[13], c34_d[13] );
  IV I21_I52 ( I21_n_0n[12], c34_d[12] );
  IV I21_I51 ( I21_n_0n[11], c34_d[11] );
  IV I21_I50 ( I21_n_0n[10], c34_d[10] );
  IV I21_I49 ( I21_n_0n[9], c34_d[9] );
  IV I21_I48 ( I21_n_0n[8], c34_d[8] );
  IV I21_I47 ( I21_n_0n[7], c34_d[7] );
  IV I21_I46 ( I21_n_0n[6], c34_d[6] );
  IV I21_I45 ( I21_n_0n[5], c34_d[5] );
  IV I21_I44 ( I21_n_0n[4], c34_d[4] );
  IV I21_I43 ( I21_n_0n[3], c34_d[3] );
  IV I21_I42 ( I21_n_0n[2], c34_d[2] );
  IV I21_I41 ( I21_n_0n[1], c34_d[1] );
  IV I21_I40 ( I21_n_0n[0], c34_d[0] );
  IV I21_I39 ( I21_nStart_0n, I21_start_0n );
  AN4 I21_I4 ( c18_a, I21_internal_0n[0], I21_internal_0n[1], I21_internal_0n[2], I21_internal_0n[3] );
  NR4 I21_I3 ( I21_internal_0n[3], I21_nCv_0n_13_, I21_nCv_0n_14_, I21_nCv_0n_15_, I21_nCv_0n_16_ );
  NR4 I21_I2 ( I21_internal_0n[2], I21_nCv_0n_9_, I21_nCv_0n_10_, I21_nCv_0n_11_, I21_nCv_0n_12_ );
  NR4 I21_I1 ( I21_internal_0n[1], I21_nCv_0n_5_, I21_nCv_0n_6_, I21_nCv_0n_7_, I21_nCv_0n_8_ );
  NR4 I21_I0 ( I21_internal_0n[0], I21_nCv_0n_1_, I21_nCv_0n_2_, I21_nCv_0n_3_, I21_nCv_0n_4_ );
  VCC I21_vcc_cell_instance ( I21_vcc );
  C2 I26_I73 ( I26_start_0n, c12_r, c12_r );
  IV I26_I55 ( I26_n_0n[15], z_0d[15] );
  IV I26_I54 ( I26_n_0n[14], z_0d[14] );
  IV I26_I53 ( I26_n_0n[13], z_0d[13] );
  IV I26_I52 ( I26_n_0n[12], z_0d[12] );
  IV I26_I51 ( I26_n_0n[11], z_0d[11] );
  IV I26_I50 ( I26_n_0n[10], z_0d[10] );
  IV I26_I49 ( I26_n_0n[9], z_0d[9] );
  IV I26_I48 ( I26_n_0n[8], z_0d[8] );
  IV I26_I47 ( I26_n_0n[7], z_0d[7] );
  IV I26_I46 ( I26_n_0n[6], z_0d[6] );
  IV I26_I45 ( I26_n_0n[5], z_0d[5] );
  IV I26_I44 ( I26_n_0n[4], z_0d[4] );
  IV I26_I43 ( I26_n_0n[3], z_0d[3] );
  IV I26_I42 ( I26_n_0n[2], z_0d[2] );
  IV I26_I41 ( I26_n_0n[1], z_0d[1] );
  IV I26_I40 ( I26_n_0n[0], z_0d[0] );
  IV I26_I39 ( I26_nStart_0n, I26_start_0n );
  AN4 I26_I4 ( c9_a, I26_internal_0n[0], I26_internal_0n[1], I26_internal_0n[2], I26_internal_0n[3] );
  NR4 I26_I3 ( I26_internal_0n[3], I26_nCv_0n_13_, I26_nCv_0n_14_, I26_nCv_0n_15_, I26_nCv_0n_16_ );
  NR4 I26_I2 ( I26_internal_0n[2], I26_nCv_0n_9_, I26_nCv_0n_10_, I26_nCv_0n_11_, I26_nCv_0n_12_ );
  NR4 I26_I1 ( I26_internal_0n[1], I26_nCv_0n_5_, I26_nCv_0n_6_, I26_nCv_0n_7_, I26_nCv_0n_8_ );
  NR4 I26_I0 ( I26_internal_0n[0], I26_nCv_0n_1_, I26_nCv_0n_2_, I26_nCv_0n_3_, I26_nCv_0n_4_ );
  VCC I26_vcc_cell_instance ( I26_vcc );
  EO I16_I13_I5 ( I16_addOut_0n_0_, I16_I13_ha, I16_vcc );
  EO I16_I13_I4 ( I16_I13_ha, I16_n_0n[0], z_0d[0] );
  NR2 I16_I13_I1 ( I16_I13_cv, I16_nStart_0n, I16_nStart_0n );
  IV I16_I13_I0 ( I16_I13_start, I16_nStart_0n );
  EO I16_I14_I5 ( I16_addOut_0n_1_, I16_I14_ha, I16_c_0n_1_ );
  EO I16_I14_I4 ( I16_I14_ha, I16_n_0n[1], z_0d[1] );
  NR2 I16_I14_I1 ( I16_I14_cv, I16_nStart_0n, I16_nCv_0n_1_ );
  IV I16_I14_I0 ( I16_I14_start, I16_nStart_0n );
  EO I16_I15_I5 ( I16_addOut_0n_2_, I16_I15_ha, I16_c_0n_2_ );
  EO I16_I15_I4 ( I16_I15_ha, I16_n_0n[2], z_0d[2] );
  NR2 I16_I15_I1 ( I16_I15_cv, I16_nStart_0n, I16_nCv_0n_2_ );
  IV I16_I15_I0 ( I16_I15_start, I16_nStart_0n );
  EO I16_I16_I5 ( I16_addOut_0n_3_, I16_I16_ha, I16_c_0n_3_ );
  EO I16_I16_I4 ( I16_I16_ha, I16_n_0n[3], z_0d[3] );
  NR2 I16_I16_I1 ( I16_I16_cv, I16_nStart_0n, I16_nCv_0n_3_ );
  IV I16_I16_I0 ( I16_I16_start, I16_nStart_0n );
  EO I16_I17_I5 ( I16_addOut_0n_4_, I16_I17_ha, I16_c_0n_4_ );
  EO I16_I17_I4 ( I16_I17_ha, I16_n_0n[4], z_0d[4] );
  NR2 I16_I17_I1 ( I16_I17_cv, I16_nStart_0n, I16_nCv_0n_4_ );
  IV I16_I17_I0 ( I16_I17_start, I16_nStart_0n );
  EO I16_I18_I5 ( I16_addOut_0n_5_, I16_I18_ha, I16_c_0n_5_ );
  EO I16_I18_I4 ( I16_I18_ha, I16_n_0n[5], z_0d[5] );
  NR2 I16_I18_I1 ( I16_I18_cv, I16_nStart_0n, I16_nCv_0n_5_ );
  IV I16_I18_I0 ( I16_I18_start, I16_nStart_0n );
  EO I16_I19_I5 ( I16_addOut_0n_6_, I16_I19_ha, I16_c_0n_6_ );
  EO I16_I19_I4 ( I16_I19_ha, I16_n_0n[6], z_0d[6] );
  NR2 I16_I19_I1 ( I16_I19_cv, I16_nStart_0n, I16_nCv_0n_6_ );
  IV I16_I19_I0 ( I16_I19_start, I16_nStart_0n );
  EO I16_I20_I5 ( I16_addOut_0n_7_, I16_I20_ha, I16_c_0n_7_ );
  EO I16_I20_I4 ( I16_I20_ha, I16_n_0n[7], z_0d[7] );
  NR2 I16_I20_I1 ( I16_I20_cv, I16_nStart_0n, I16_nCv_0n_7_ );
  IV I16_I20_I0 ( I16_I20_start, I16_nStart_0n );
  EO I16_I21_I5 ( I16_addOut_0n_8_, I16_I21_ha, I16_c_0n_8_ );
  EO I16_I21_I4 ( I16_I21_ha, I16_n_0n[8], z_0d[8] );
  NR2 I16_I21_I1 ( I16_I21_cv, I16_nStart_0n, I16_nCv_0n_8_ );
  IV I16_I21_I0 ( I16_I21_start, I16_nStart_0n );
  EO I16_I22_I5 ( I16_addOut_0n_9_, I16_I22_ha, I16_c_0n_9_ );
  EO I16_I22_I4 ( I16_I22_ha, I16_n_0n[9], z_0d[9] );
  NR2 I16_I22_I1 ( I16_I22_cv, I16_nStart_0n, I16_nCv_0n_9_ );
  IV I16_I22_I0 ( I16_I22_start, I16_nStart_0n );
  EO I16_I23_I5 ( I16_addOut_0n_10_, I16_I23_ha, I16_c_0n_10_ );
  EO I16_I23_I4 ( I16_I23_ha, I16_n_0n[10], z_0d[10] );
  NR2 I16_I23_I1 ( I16_I23_cv, I16_nStart_0n, I16_nCv_0n_10_ );
  IV I16_I23_I0 ( I16_I23_start, I16_nStart_0n );
  EO I16_I24_I5 ( I16_addOut_0n_11_, I16_I24_ha, I16_c_0n_11_ );
  EO I16_I24_I4 ( I16_I24_ha, I16_n_0n[11], z_0d[11] );
  NR2 I16_I24_I1 ( I16_I24_cv, I16_nStart_0n, I16_nCv_0n_11_ );
  IV I16_I24_I0 ( I16_I24_start, I16_nStart_0n );
  EO I16_I25_I5 ( I16_addOut_0n_12_, I16_I25_ha, I16_c_0n_12_ );
  EO I16_I25_I4 ( I16_I25_ha, I16_n_0n[12], z_0d[12] );
  NR2 I16_I25_I1 ( I16_I25_cv, I16_nStart_0n, I16_nCv_0n_12_ );
  IV I16_I25_I0 ( I16_I25_start, I16_nStart_0n );
  EO I16_I26_I5 ( I16_addOut_0n_13_, I16_I26_ha, I16_c_0n_13_ );
  EO I16_I26_I4 ( I16_I26_ha, I16_n_0n[13], z_0d[13] );
  NR2 I16_I26_I1 ( I16_I26_cv, I16_nStart_0n, I16_nCv_0n_13_ );
  IV I16_I26_I0 ( I16_I26_start, I16_nStart_0n );
  EO I16_I27_I5 ( I16_addOut_0n_14_, I16_I27_ha, I16_c_0n_14_ );
  EO I16_I27_I4 ( I16_I27_ha, I16_n_0n[14], z_0d[14] );
  NR2 I16_I27_I1 ( I16_I27_cv, I16_nStart_0n, I16_nCv_0n_14_ );
  IV I16_I27_I0 ( I16_I27_start, I16_nStart_0n );
  EO I16_I28_I5 ( I16_addOut_0n_15_, I16_I28_ha, I16_c_0n_15_ );
  EO I16_I28_I4 ( I16_I28_ha, I16_n_0n[15], z_0d[15] );
  NR2 I16_I28_I1 ( I16_I28_cv, I16_nStart_0n, I16_nCv_0n_15_ );
  IV I16_I28_I0 ( I16_I28_start, I16_nStart_0n );
  EO I21_I21_I5 ( c18_d[0], I21_I21_ha, I21_vcc );
  EO I21_I21_I4 ( I21_I21_ha, I21_n_0n[0], z_0d[0] );
  NR2 I21_I21_I1 ( I21_I21_cv, I21_nStart_0n, I21_nStart_0n );
  IV I21_I21_I0 ( I21_I21_start, I21_nStart_0n );
  EO I21_I22_I5 ( c18_d[1], I21_I22_ha, I21_c_0n[1] );
  EO I21_I22_I4 ( I21_I22_ha, I21_n_0n[1], z_0d[1] );
  NR2 I21_I22_I1 ( I21_I22_cv, I21_nStart_0n, I21_nCv_0n_1_ );
  IV I21_I22_I0 ( I21_I22_start, I21_nStart_0n );
  EO I21_I23_I5 ( c18_d[2], I21_I23_ha, I21_c_0n[2] );
  EO I21_I23_I4 ( I21_I23_ha, I21_n_0n[2], z_0d[2] );
  NR2 I21_I23_I1 ( I21_I23_cv, I21_nStart_0n, I21_nCv_0n_2_ );
  IV I21_I23_I0 ( I21_I23_start, I21_nStart_0n );
  EO I21_I24_I5 ( c18_d[3], I21_I24_ha, I21_c_0n[3] );
  EO I21_I24_I4 ( I21_I24_ha, I21_n_0n[3], z_0d[3] );
  NR2 I21_I24_I1 ( I21_I24_cv, I21_nStart_0n, I21_nCv_0n_3_ );
  IV I21_I24_I0 ( I21_I24_start, I21_nStart_0n );
  EO I21_I25_I5 ( c18_d[4], I21_I25_ha, I21_c_0n[4] );
  EO I21_I25_I4 ( I21_I25_ha, I21_n_0n[4], z_0d[4] );
  NR2 I21_I25_I1 ( I21_I25_cv, I21_nStart_0n, I21_nCv_0n_4_ );
  IV I21_I25_I0 ( I21_I25_start, I21_nStart_0n );
  EO I21_I26_I5 ( c18_d[5], I21_I26_ha, I21_c_0n[5] );
  EO I21_I26_I4 ( I21_I26_ha, I21_n_0n[5], z_0d[5] );
  NR2 I21_I26_I1 ( I21_I26_cv, I21_nStart_0n, I21_nCv_0n_5_ );
  IV I21_I26_I0 ( I21_I26_start, I21_nStart_0n );
  EO I21_I27_I5 ( c18_d[6], I21_I27_ha, I21_c_0n[6] );
  EO I21_I27_I4 ( I21_I27_ha, I21_n_0n[6], z_0d[6] );
  NR2 I21_I27_I1 ( I21_I27_cv, I21_nStart_0n, I21_nCv_0n_6_ );
  IV I21_I27_I0 ( I21_I27_start, I21_nStart_0n );
  EO I21_I28_I5 ( c18_d[7], I21_I28_ha, I21_c_0n[7] );
  EO I21_I28_I4 ( I21_I28_ha, I21_n_0n[7], z_0d[7] );
  NR2 I21_I28_I1 ( I21_I28_cv, I21_nStart_0n, I21_nCv_0n_7_ );
  IV I21_I28_I0 ( I21_I28_start, I21_nStart_0n );
  EO I21_I29_I5 ( c18_d[8], I21_I29_ha, I21_c_0n[8] );
  EO I21_I29_I4 ( I21_I29_ha, I21_n_0n[8], z_0d[8] );
  NR2 I21_I29_I1 ( I21_I29_cv, I21_nStart_0n, I21_nCv_0n_8_ );
  IV I21_I29_I0 ( I21_I29_start, I21_nStart_0n );
  EO I21_I30_I5 ( c18_d[9], I21_I30_ha, I21_c_0n[9] );
  EO I21_I30_I4 ( I21_I30_ha, I21_n_0n[9], z_0d[9] );
  NR2 I21_I30_I1 ( I21_I30_cv, I21_nStart_0n, I21_nCv_0n_9_ );
  IV I21_I30_I0 ( I21_I30_start, I21_nStart_0n );
  EO I21_I31_I5 ( c18_d[10], I21_I31_ha, I21_c_0n[10] );
  EO I21_I31_I4 ( I21_I31_ha, I21_n_0n[10], z_0d[10] );
  NR2 I21_I31_I1 ( I21_I31_cv, I21_nStart_0n, I21_nCv_0n_10_ );
  IV I21_I31_I0 ( I21_I31_start, I21_nStart_0n );
  EO I21_I32_I5 ( c18_d[11], I21_I32_ha, I21_c_0n[11] );
  EO I21_I32_I4 ( I21_I32_ha, I21_n_0n[11], z_0d[11] );
  NR2 I21_I32_I1 ( I21_I32_cv, I21_nStart_0n, I21_nCv_0n_11_ );
  IV I21_I32_I0 ( I21_I32_start, I21_nStart_0n );
  EO I21_I33_I5 ( c18_d[12], I21_I33_ha, I21_c_0n[12] );
  EO I21_I33_I4 ( I21_I33_ha, I21_n_0n[12], z_0d[12] );
  NR2 I21_I33_I1 ( I21_I33_cv, I21_nStart_0n, I21_nCv_0n_12_ );
  IV I21_I33_I0 ( I21_I33_start, I21_nStart_0n );
  EO I21_I34_I5 ( c18_d[13], I21_I34_ha, I21_c_0n[13] );
  EO I21_I34_I4 ( I21_I34_ha, I21_n_0n[13], z_0d[13] );
  NR2 I21_I34_I1 ( I21_I34_cv, I21_nStart_0n, I21_nCv_0n_13_ );
  IV I21_I34_I0 ( I21_I34_start, I21_nStart_0n );
  EO I21_I35_I5 ( c18_d[14], I21_I35_ha, I21_c_0n[14] );
  EO I21_I35_I4 ( I21_I35_ha, I21_n_0n[14], z_0d[14] );
  NR2 I21_I35_I1 ( I21_I35_cv, I21_nStart_0n, I21_nCv_0n_14_ );
  IV I21_I35_I0 ( I21_I35_start, I21_nStart_0n );
  EO I21_I36_I5 ( c18_d[15], I21_I36_ha, I21_c_0n[15] );
  EO I21_I36_I4 ( I21_I36_ha, I21_n_0n[15], z_0d[15] );
  NR2 I21_I36_I1 ( I21_I36_cv, I21_nStart_0n, I21_nCv_0n_15_ );
  IV I21_I36_I0 ( I21_I36_start, I21_nStart_0n );
  EO I26_I21_I5 ( c9_d[0], I26_I21_ha, I26_vcc );
  EO I26_I21_I4 ( I26_I21_ha, I26_n_0n[0], c34_d[0] );
  NR2 I26_I21_I1 ( I26_I21_cv, I26_nStart_0n, I26_nStart_0n );
  IV I26_I21_I0 ( I26_I21_start, I26_nStart_0n );
  EO I26_I22_I5 ( c9_d[1], I26_I22_ha, I26_c_0n[1] );
  EO I26_I22_I4 ( I26_I22_ha, I26_n_0n[1], c34_d[1] );
  NR2 I26_I22_I1 ( I26_I22_cv, I26_nStart_0n, I26_nCv_0n_1_ );
  IV I26_I22_I0 ( I26_I22_start, I26_nStart_0n );
  EO I26_I23_I5 ( c9_d[2], I26_I23_ha, I26_c_0n[2] );
  EO I26_I23_I4 ( I26_I23_ha, I26_n_0n[2], c34_d[2] );
  NR2 I26_I23_I1 ( I26_I23_cv, I26_nStart_0n, I26_nCv_0n_2_ );
  IV I26_I23_I0 ( I26_I23_start, I26_nStart_0n );
  EO I26_I24_I5 ( c9_d[3], I26_I24_ha, I26_c_0n[3] );
  EO I26_I24_I4 ( I26_I24_ha, I26_n_0n[3], c34_d[3] );
  NR2 I26_I24_I1 ( I26_I24_cv, I26_nStart_0n, I26_nCv_0n_3_ );
  IV I26_I24_I0 ( I26_I24_start, I26_nStart_0n );
  EO I26_I25_I5 ( c9_d[4], I26_I25_ha, I26_c_0n[4] );
  EO I26_I25_I4 ( I26_I25_ha, I26_n_0n[4], c34_d[4] );
  NR2 I26_I25_I1 ( I26_I25_cv, I26_nStart_0n, I26_nCv_0n_4_ );
  IV I26_I25_I0 ( I26_I25_start, I26_nStart_0n );
  EO I26_I26_I5 ( c9_d[5], I26_I26_ha, I26_c_0n[5] );
  EO I26_I26_I4 ( I26_I26_ha, I26_n_0n[5], c34_d[5] );
  NR2 I26_I26_I1 ( I26_I26_cv, I26_nStart_0n, I26_nCv_0n_5_ );
  IV I26_I26_I0 ( I26_I26_start, I26_nStart_0n );
  EO I26_I27_I5 ( c9_d[6], I26_I27_ha, I26_c_0n[6] );
  EO I26_I27_I4 ( I26_I27_ha, I26_n_0n[6], c34_d[6] );
  NR2 I26_I27_I1 ( I26_I27_cv, I26_nStart_0n, I26_nCv_0n_6_ );
  IV I26_I27_I0 ( I26_I27_start, I26_nStart_0n );
  EO I26_I28_I5 ( c9_d[7], I26_I28_ha, I26_c_0n[7] );
  EO I26_I28_I4 ( I26_I28_ha, I26_n_0n[7], c34_d[7] );
  NR2 I26_I28_I1 ( I26_I28_cv, I26_nStart_0n, I26_nCv_0n_7_ );
  IV I26_I28_I0 ( I26_I28_start, I26_nStart_0n );
  EO I26_I29_I5 ( c9_d[8], I26_I29_ha, I26_c_0n[8] );
  EO I26_I29_I4 ( I26_I29_ha, I26_n_0n[8], c34_d[8] );
  NR2 I26_I29_I1 ( I26_I29_cv, I26_nStart_0n, I26_nCv_0n_8_ );
  IV I26_I29_I0 ( I26_I29_start, I26_nStart_0n );
  EO I26_I30_I5 ( c9_d[9], I26_I30_ha, I26_c_0n[9] );
  EO I26_I30_I4 ( I26_I30_ha, I26_n_0n[9], c34_d[9] );
  NR2 I26_I30_I1 ( I26_I30_cv, I26_nStart_0n, I26_nCv_0n_9_ );
  IV I26_I30_I0 ( I26_I30_start, I26_nStart_0n );
  EO I26_I31_I5 ( c9_d[10], I26_I31_ha, I26_c_0n[10] );
  EO I26_I31_I4 ( I26_I31_ha, I26_n_0n[10], c34_d[10] );
  NR2 I26_I31_I1 ( I26_I31_cv, I26_nStart_0n, I26_nCv_0n_10_ );
  IV I26_I31_I0 ( I26_I31_start, I26_nStart_0n );
  EO I26_I32_I5 ( c9_d[11], I26_I32_ha, I26_c_0n[11] );
  EO I26_I32_I4 ( I26_I32_ha, I26_n_0n[11], c34_d[11] );
  NR2 I26_I32_I1 ( I26_I32_cv, I26_nStart_0n, I26_nCv_0n_11_ );
  IV I26_I32_I0 ( I26_I32_start, I26_nStart_0n );
  EO I26_I33_I5 ( c9_d[12], I26_I33_ha, I26_c_0n[12] );
  EO I26_I33_I4 ( I26_I33_ha, I26_n_0n[12], c34_d[12] );
  NR2 I26_I33_I1 ( I26_I33_cv, I26_nStart_0n, I26_nCv_0n_12_ );
  IV I26_I33_I0 ( I26_I33_start, I26_nStart_0n );
  EO I26_I34_I5 ( c9_d[13], I26_I34_ha, I26_c_0n[13] );
  EO I26_I34_I4 ( I26_I34_ha, I26_n_0n[13], c34_d[13] );
  NR2 I26_I34_I1 ( I26_I34_cv, I26_nStart_0n, I26_nCv_0n_13_ );
  IV I26_I34_I0 ( I26_I34_start, I26_nStart_0n );
  EO I26_I35_I5 ( c9_d[14], I26_I35_ha, I26_c_0n[14] );
  EO I26_I35_I4 ( I26_I35_ha, I26_n_0n[14], c34_d[14] );
  NR2 I26_I35_I1 ( I26_I35_cv, I26_nStart_0n, I26_nCv_0n_14_ );
  IV I26_I35_I0 ( I26_I35_start, I26_nStart_0n );
  EO I26_I36_I5 ( c9_d[15], I26_I36_ha, I26_c_0n[15] );
  EO I26_I36_I4 ( I26_I36_ha, I26_n_0n[15], c34_d[15] );
  NR2 I26_I36_I1 ( I26_I36_cv, I26_nStart_0n, I26_nCv_0n_15_ );
  IV I26_I36_I0 ( I26_I36_start, I26_nStart_0n );
  IV I16_I13_I2_I1 ( I16_I13_I2_nsel_0n, I16_I13_ha );
  IV I16_I14_I2_I1 ( I16_I14_I2_nsel_0n, I16_I14_ha );
  IV I16_I15_I2_I1 ( I16_I15_I2_nsel_0n, I16_I15_ha );
  IV I16_I16_I2_I1 ( I16_I16_I2_nsel_0n, I16_I16_ha );
  IV I16_I17_I2_I1 ( I16_I17_I2_nsel_0n, I16_I17_ha );
  IV I16_I18_I2_I1 ( I16_I18_I2_nsel_0n, I16_I18_ha );
  IV I16_I19_I2_I1 ( I16_I19_I2_nsel_0n, I16_I19_ha );
  IV I16_I20_I2_I1 ( I16_I20_I2_nsel_0n, I16_I20_ha );
  IV I16_I21_I2_I1 ( I16_I21_I2_nsel_0n, I16_I21_ha );
  IV I16_I22_I2_I1 ( I16_I22_I2_nsel_0n, I16_I22_ha );
  IV I16_I23_I2_I1 ( I16_I23_I2_nsel_0n, I16_I23_ha );
  IV I16_I24_I2_I1 ( I16_I24_I2_nsel_0n, I16_I24_ha );
  IV I16_I25_I2_I1 ( I16_I25_I2_nsel_0n, I16_I25_ha );
  IV I16_I26_I2_I1 ( I16_I26_I2_nsel_0n, I16_I26_ha );
  IV I16_I27_I2_I1 ( I16_I27_I2_nsel_0n, I16_I27_ha );
  IV I16_I28_I2_I1 ( I16_I28_I2_nsel_0n, I16_I28_ha );
  IV I21_I21_I2_I1 ( I21_I21_I2_nsel_0n, I21_I21_ha );
  IV I21_I22_I2_I1 ( I21_I22_I2_nsel_0n, I21_I22_ha );
  IV I21_I23_I2_I1 ( I21_I23_I2_nsel_0n, I21_I23_ha );
  IV I21_I24_I2_I1 ( I21_I24_I2_nsel_0n, I21_I24_ha );
  IV I21_I25_I2_I1 ( I21_I25_I2_nsel_0n, I21_I25_ha );
  IV I21_I26_I2_I1 ( I21_I26_I2_nsel_0n, I21_I26_ha );
  IV I21_I27_I2_I1 ( I21_I27_I2_nsel_0n, I21_I27_ha );
  IV I21_I28_I2_I1 ( I21_I28_I2_nsel_0n, I21_I28_ha );
  IV I21_I29_I2_I1 ( I21_I29_I2_nsel_0n, I21_I29_ha );
  IV I21_I30_I2_I1 ( I21_I30_I2_nsel_0n, I21_I30_ha );
  IV I21_I31_I2_I1 ( I21_I31_I2_nsel_0n, I21_I31_ha );
  IV I21_I32_I2_I1 ( I21_I32_I2_nsel_0n, I21_I32_ha );
  IV I21_I33_I2_I1 ( I21_I33_I2_nsel_0n, I21_I33_ha );
  IV I21_I34_I2_I1 ( I21_I34_I2_nsel_0n, I21_I34_ha );
  IV I21_I35_I2_I1 ( I21_I35_I2_nsel_0n, I21_I35_ha );
  IV I21_I36_I2_I1 ( I21_I36_I2_nsel_0n, I21_I36_ha );
  IV I26_I21_I2_I1 ( I26_I21_I2_nsel_0n, I26_I21_ha );
  IV I26_I22_I2_I1 ( I26_I22_I2_nsel_0n, I26_I22_ha );
  IV I26_I23_I2_I1 ( I26_I23_I2_nsel_0n, I26_I23_ha );
  IV I26_I24_I2_I1 ( I26_I24_I2_nsel_0n, I26_I24_ha );
  IV I26_I25_I2_I1 ( I26_I25_I2_nsel_0n, I26_I25_ha );
  IV I26_I26_I2_I1 ( I26_I26_I2_nsel_0n, I26_I26_ha );
  IV I26_I27_I2_I1 ( I26_I27_I2_nsel_0n, I26_I27_ha );
  IV I26_I28_I2_I1 ( I26_I28_I2_nsel_0n, I26_I28_ha );
  IV I26_I29_I2_I1 ( I26_I29_I2_nsel_0n, I26_I29_ha );
  IV I26_I30_I2_I1 ( I26_I30_I2_nsel_0n, I26_I30_ha );
  IV I26_I31_I2_I1 ( I26_I31_I2_nsel_0n, I26_I31_ha );
  IV I26_I32_I2_I1 ( I26_I32_I2_nsel_0n, I26_I32_ha );
  IV I26_I33_I2_I1 ( I26_I33_I2_nsel_0n, I26_I33_ha );
  IV I26_I34_I2_I1 ( I26_I34_I2_nsel_0n, I26_I34_ha );
  IV I26_I35_I2_I1 ( I26_I35_I2_nsel_0n, I26_I35_ha );
  IV I26_I36_I2_I1 ( I26_I36_I2_nsel_0n, I26_I36_ha );
  AN2 I16_I13_I2_I0_I2 ( I16_I13_I2_I0_int_0n[0], I16_I13_start, I16_I13_I2_nsel_0n );
  AN2 I16_I13_I2_I0_I1 ( I16_I13_I2_I0_int_0n[1], I16_I13_cv, I16_I13_ha );
  NR2 I16_I13_I2_I0_I0 ( I16_nCv_0n_1_, I16_I13_I2_I0_int_0n[0], I16_I13_I2_I0_int_0n[1] );
  AN2 I16_I14_I2_I0_I2 ( I16_I14_I2_I0_int_0n[0], I16_I14_start, I16_I14_I2_nsel_0n );
  AN2 I16_I14_I2_I0_I1 ( I16_I14_I2_I0_int_0n[1], I16_I14_cv, I16_I14_ha );
  NR2 I16_I14_I2_I0_I0 ( I16_nCv_0n_2_, I16_I14_I2_I0_int_0n[0], I16_I14_I2_I0_int_0n[1] );
  AN2 I16_I15_I2_I0_I2 ( I16_I15_I2_I0_int_0n[0], I16_I15_start, I16_I15_I2_nsel_0n );
  AN2 I16_I15_I2_I0_I1 ( I16_I15_I2_I0_int_0n[1], I16_I15_cv, I16_I15_ha );
  NR2 I16_I15_I2_I0_I0 ( I16_nCv_0n_3_, I16_I15_I2_I0_int_0n[0], I16_I15_I2_I0_int_0n[1] );
  AN2 I16_I16_I2_I0_I2 ( I16_I16_I2_I0_int_0n[0], I16_I16_start, I16_I16_I2_nsel_0n );
  AN2 I16_I16_I2_I0_I1 ( I16_I16_I2_I0_int_0n[1], I16_I16_cv, I16_I16_ha );
  NR2 I16_I16_I2_I0_I0 ( I16_nCv_0n_4_, I16_I16_I2_I0_int_0n[0], I16_I16_I2_I0_int_0n[1] );
  AN2 I16_I17_I2_I0_I2 ( I16_I17_I2_I0_int_0n[0], I16_I17_start, I16_I17_I2_nsel_0n );
  AN2 I16_I17_I2_I0_I1 ( I16_I17_I2_I0_int_0n[1], I16_I17_cv, I16_I17_ha );
  NR2 I16_I17_I2_I0_I0 ( I16_nCv_0n_5_, I16_I17_I2_I0_int_0n[0], I16_I17_I2_I0_int_0n[1] );
  AN2 I16_I18_I2_I0_I2 ( I16_I18_I2_I0_int_0n[0], I16_I18_start, I16_I18_I2_nsel_0n );
  AN2 I16_I18_I2_I0_I1 ( I16_I18_I2_I0_int_0n[1], I16_I18_cv, I16_I18_ha );
  NR2 I16_I18_I2_I0_I0 ( I16_nCv_0n_6_, I16_I18_I2_I0_int_0n[0], I16_I18_I2_I0_int_0n[1] );
  AN2 I16_I19_I2_I0_I2 ( I16_I19_I2_I0_int_0n[0], I16_I19_start, I16_I19_I2_nsel_0n );
  AN2 I16_I19_I2_I0_I1 ( I16_I19_I2_I0_int_0n[1], I16_I19_cv, I16_I19_ha );
  NR2 I16_I19_I2_I0_I0 ( I16_nCv_0n_7_, I16_I19_I2_I0_int_0n[0], I16_I19_I2_I0_int_0n[1] );
  AN2 I16_I20_I2_I0_I2 ( I16_I20_I2_I0_int_0n[0], I16_I20_start, I16_I20_I2_nsel_0n );
  AN2 I16_I20_I2_I0_I1 ( I16_I20_I2_I0_int_0n[1], I16_I20_cv, I16_I20_ha );
  NR2 I16_I20_I2_I0_I0 ( I16_nCv_0n_8_, I16_I20_I2_I0_int_0n[0], I16_I20_I2_I0_int_0n[1] );
  AN2 I16_I21_I2_I0_I2 ( I16_I21_I2_I0_int_0n[0], I16_I21_start, I16_I21_I2_nsel_0n );
  AN2 I16_I21_I2_I0_I1 ( I16_I21_I2_I0_int_0n[1], I16_I21_cv, I16_I21_ha );
  NR2 I16_I21_I2_I0_I0 ( I16_nCv_0n_9_, I16_I21_I2_I0_int_0n[0], I16_I21_I2_I0_int_0n[1] );
  AN2 I16_I22_I2_I0_I2 ( I16_I22_I2_I0_int_0n[0], I16_I22_start, I16_I22_I2_nsel_0n );
  AN2 I16_I22_I2_I0_I1 ( I16_I22_I2_I0_int_0n[1], I16_I22_cv, I16_I22_ha );
  NR2 I16_I22_I2_I0_I0 ( I16_nCv_0n_10_, I16_I22_I2_I0_int_0n[0], I16_I22_I2_I0_int_0n[1] );
  AN2 I16_I23_I2_I0_I2 ( I16_I23_I2_I0_int_0n[0], I16_I23_start, I16_I23_I2_nsel_0n );
  AN2 I16_I23_I2_I0_I1 ( I16_I23_I2_I0_int_0n[1], I16_I23_cv, I16_I23_ha );
  NR2 I16_I23_I2_I0_I0 ( I16_nCv_0n_11_, I16_I23_I2_I0_int_0n[0], I16_I23_I2_I0_int_0n[1] );
  AN2 I16_I24_I2_I0_I2 ( I16_I24_I2_I0_int_0n[0], I16_I24_start, I16_I24_I2_nsel_0n );
  AN2 I16_I24_I2_I0_I1 ( I16_I24_I2_I0_int_0n[1], I16_I24_cv, I16_I24_ha );
  NR2 I16_I24_I2_I0_I0 ( I16_nCv_0n_12_, I16_I24_I2_I0_int_0n[0], I16_I24_I2_I0_int_0n[1] );
  AN2 I16_I25_I2_I0_I2 ( I16_I25_I2_I0_int_0n[0], I16_I25_start, I16_I25_I2_nsel_0n );
  AN2 I16_I25_I2_I0_I1 ( I16_I25_I2_I0_int_0n[1], I16_I25_cv, I16_I25_ha );
  NR2 I16_I25_I2_I0_I0 ( I16_nCv_0n_13_, I16_I25_I2_I0_int_0n[0], I16_I25_I2_I0_int_0n[1] );
  AN2 I16_I26_I2_I0_I2 ( I16_I26_I2_I0_int_0n[0], I16_I26_start, I16_I26_I2_nsel_0n );
  AN2 I16_I26_I2_I0_I1 ( I16_I26_I2_I0_int_0n[1], I16_I26_cv, I16_I26_ha );
  NR2 I16_I26_I2_I0_I0 ( I16_nCv_0n_14_, I16_I26_I2_I0_int_0n[0], I16_I26_I2_I0_int_0n[1] );
  AN2 I16_I27_I2_I0_I2 ( I16_I27_I2_I0_int_0n[0], I16_I27_start, I16_I27_I2_nsel_0n );
  AN2 I16_I27_I2_I0_I1 ( I16_I27_I2_I0_int_0n[1], I16_I27_cv, I16_I27_ha );
  NR2 I16_I27_I2_I0_I0 ( I16_nCv_0n_15_, I16_I27_I2_I0_int_0n[0], I16_I27_I2_I0_int_0n[1] );
  AN2 I16_I28_I2_I0_I2 ( I16_I28_I2_I0_int_0n[0], I16_I28_start, I16_I28_I2_nsel_0n );
  AN2 I16_I28_I2_I0_I1 ( I16_I28_I2_I0_int_0n[1], I16_I28_cv, I16_I28_ha );
  NR2 I16_I28_I2_I0_I0 ( I16_nCv_0n_16_, I16_I28_I2_I0_int_0n[0], I16_I28_I2_I0_int_0n[1] );
  AN2 I21_I21_I2_I0_I2 ( I21_I21_I2_I0_int_0n[0], I21_I21_start, I21_I21_I2_nsel_0n );
  AN2 I21_I21_I2_I0_I1 ( I21_I21_I2_I0_int_0n[1], I21_I21_cv, I21_I21_ha );
  NR2 I21_I21_I2_I0_I0 ( I21_nCv_0n_1_, I21_I21_I2_I0_int_0n[0], I21_I21_I2_I0_int_0n[1] );
  AN2 I21_I22_I2_I0_I2 ( I21_I22_I2_I0_int_0n[0], I21_I22_start, I21_I22_I2_nsel_0n );
  AN2 I21_I22_I2_I0_I1 ( I21_I22_I2_I0_int_0n[1], I21_I22_cv, I21_I22_ha );
  NR2 I21_I22_I2_I0_I0 ( I21_nCv_0n_2_, I21_I22_I2_I0_int_0n[0], I21_I22_I2_I0_int_0n[1] );
  AN2 I21_I23_I2_I0_I2 ( I21_I23_I2_I0_int_0n[0], I21_I23_start, I21_I23_I2_nsel_0n );
  AN2 I21_I23_I2_I0_I1 ( I21_I23_I2_I0_int_0n[1], I21_I23_cv, I21_I23_ha );
  NR2 I21_I23_I2_I0_I0 ( I21_nCv_0n_3_, I21_I23_I2_I0_int_0n[0], I21_I23_I2_I0_int_0n[1] );
  AN2 I21_I24_I2_I0_I2 ( I21_I24_I2_I0_int_0n[0], I21_I24_start, I21_I24_I2_nsel_0n );
  AN2 I21_I24_I2_I0_I1 ( I21_I24_I2_I0_int_0n[1], I21_I24_cv, I21_I24_ha );
  NR2 I21_I24_I2_I0_I0 ( I21_nCv_0n_4_, I21_I24_I2_I0_int_0n[0], I21_I24_I2_I0_int_0n[1] );
  AN2 I21_I25_I2_I0_I2 ( I21_I25_I2_I0_int_0n[0], I21_I25_start, I21_I25_I2_nsel_0n );
  AN2 I21_I25_I2_I0_I1 ( I21_I25_I2_I0_int_0n[1], I21_I25_cv, I21_I25_ha );
  NR2 I21_I25_I2_I0_I0 ( I21_nCv_0n_5_, I21_I25_I2_I0_int_0n[0], I21_I25_I2_I0_int_0n[1] );
  AN2 I21_I26_I2_I0_I2 ( I21_I26_I2_I0_int_0n[0], I21_I26_start, I21_I26_I2_nsel_0n );
  AN2 I21_I26_I2_I0_I1 ( I21_I26_I2_I0_int_0n[1], I21_I26_cv, I21_I26_ha );
  NR2 I21_I26_I2_I0_I0 ( I21_nCv_0n_6_, I21_I26_I2_I0_int_0n[0], I21_I26_I2_I0_int_0n[1] );
  AN2 I21_I27_I2_I0_I2 ( I21_I27_I2_I0_int_0n[0], I21_I27_start, I21_I27_I2_nsel_0n );
  AN2 I21_I27_I2_I0_I1 ( I21_I27_I2_I0_int_0n[1], I21_I27_cv, I21_I27_ha );
  NR2 I21_I27_I2_I0_I0 ( I21_nCv_0n_7_, I21_I27_I2_I0_int_0n[0], I21_I27_I2_I0_int_0n[1] );
  AN2 I21_I28_I2_I0_I2 ( I21_I28_I2_I0_int_0n[0], I21_I28_start, I21_I28_I2_nsel_0n );
  AN2 I21_I28_I2_I0_I1 ( I21_I28_I2_I0_int_0n[1], I21_I28_cv, I21_I28_ha );
  NR2 I21_I28_I2_I0_I0 ( I21_nCv_0n_8_, I21_I28_I2_I0_int_0n[0], I21_I28_I2_I0_int_0n[1] );
  AN2 I21_I29_I2_I0_I2 ( I21_I29_I2_I0_int_0n[0], I21_I29_start, I21_I29_I2_nsel_0n );
  AN2 I21_I29_I2_I0_I1 ( I21_I29_I2_I0_int_0n[1], I21_I29_cv, I21_I29_ha );
  NR2 I21_I29_I2_I0_I0 ( I21_nCv_0n_9_, I21_I29_I2_I0_int_0n[0], I21_I29_I2_I0_int_0n[1] );
  AN2 I21_I30_I2_I0_I2 ( I21_I30_I2_I0_int_0n[0], I21_I30_start, I21_I30_I2_nsel_0n );
  AN2 I21_I30_I2_I0_I1 ( I21_I30_I2_I0_int_0n[1], I21_I30_cv, I21_I30_ha );
  NR2 I21_I30_I2_I0_I0 ( I21_nCv_0n_10_, I21_I30_I2_I0_int_0n[0], I21_I30_I2_I0_int_0n[1] );
  AN2 I21_I31_I2_I0_I2 ( I21_I31_I2_I0_int_0n[0], I21_I31_start, I21_I31_I2_nsel_0n );
  AN2 I21_I31_I2_I0_I1 ( I21_I31_I2_I0_int_0n[1], I21_I31_cv, I21_I31_ha );
  NR2 I21_I31_I2_I0_I0 ( I21_nCv_0n_11_, I21_I31_I2_I0_int_0n[0], I21_I31_I2_I0_int_0n[1] );
  AN2 I21_I32_I2_I0_I2 ( I21_I32_I2_I0_int_0n[0], I21_I32_start, I21_I32_I2_nsel_0n );
  AN2 I21_I32_I2_I0_I1 ( I21_I32_I2_I0_int_0n[1], I21_I32_cv, I21_I32_ha );
  NR2 I21_I32_I2_I0_I0 ( I21_nCv_0n_12_, I21_I32_I2_I0_int_0n[0], I21_I32_I2_I0_int_0n[1] );
  AN2 I21_I33_I2_I0_I2 ( I21_I33_I2_I0_int_0n[0], I21_I33_start, I21_I33_I2_nsel_0n );
  AN2 I21_I33_I2_I0_I1 ( I21_I33_I2_I0_int_0n[1], I21_I33_cv, I21_I33_ha );
  NR2 I21_I33_I2_I0_I0 ( I21_nCv_0n_13_, I21_I33_I2_I0_int_0n[0], I21_I33_I2_I0_int_0n[1] );
  AN2 I21_I34_I2_I0_I2 ( I21_I34_I2_I0_int_0n[0], I21_I34_start, I21_I34_I2_nsel_0n );
  AN2 I21_I34_I2_I0_I1 ( I21_I34_I2_I0_int_0n[1], I21_I34_cv, I21_I34_ha );
  NR2 I21_I34_I2_I0_I0 ( I21_nCv_0n_14_, I21_I34_I2_I0_int_0n[0], I21_I34_I2_I0_int_0n[1] );
  AN2 I21_I35_I2_I0_I2 ( I21_I35_I2_I0_int_0n[0], I21_I35_start, I21_I35_I2_nsel_0n );
  AN2 I21_I35_I2_I0_I1 ( I21_I35_I2_I0_int_0n[1], I21_I35_cv, I21_I35_ha );
  NR2 I21_I35_I2_I0_I0 ( I21_nCv_0n_15_, I21_I35_I2_I0_int_0n[0], I21_I35_I2_I0_int_0n[1] );
  AN2 I21_I36_I2_I0_I2 ( I21_I36_I2_I0_int_0n[0], I21_I36_start, I21_I36_I2_nsel_0n );
  AN2 I21_I36_I2_I0_I1 ( I21_I36_I2_I0_int_0n[1], I21_I36_cv, I21_I36_ha );
  NR2 I21_I36_I2_I0_I0 ( I21_nCv_0n_16_, I21_I36_I2_I0_int_0n[0], I21_I36_I2_I0_int_0n[1] );
  AN2 I26_I21_I2_I0_I2 ( I26_I21_I2_I0_int_0n[0], I26_I21_start, I26_I21_I2_nsel_0n );
  AN2 I26_I21_I2_I0_I1 ( I26_I21_I2_I0_int_0n[1], I26_I21_cv, I26_I21_ha );
  NR2 I26_I21_I2_I0_I0 ( I26_nCv_0n_1_, I26_I21_I2_I0_int_0n[0], I26_I21_I2_I0_int_0n[1] );
  AN2 I26_I22_I2_I0_I2 ( I26_I22_I2_I0_int_0n[0], I26_I22_start, I26_I22_I2_nsel_0n );
  AN2 I26_I22_I2_I0_I1 ( I26_I22_I2_I0_int_0n[1], I26_I22_cv, I26_I22_ha );
  NR2 I26_I22_I2_I0_I0 ( I26_nCv_0n_2_, I26_I22_I2_I0_int_0n[0], I26_I22_I2_I0_int_0n[1] );
  AN2 I26_I23_I2_I0_I2 ( I26_I23_I2_I0_int_0n[0], I26_I23_start, I26_I23_I2_nsel_0n );
  AN2 I26_I23_I2_I0_I1 ( I26_I23_I2_I0_int_0n[1], I26_I23_cv, I26_I23_ha );
  NR2 I26_I23_I2_I0_I0 ( I26_nCv_0n_3_, I26_I23_I2_I0_int_0n[0], I26_I23_I2_I0_int_0n[1] );
  AN2 I26_I24_I2_I0_I2 ( I26_I24_I2_I0_int_0n[0], I26_I24_start, I26_I24_I2_nsel_0n );
  AN2 I26_I24_I2_I0_I1 ( I26_I24_I2_I0_int_0n[1], I26_I24_cv, I26_I24_ha );
  NR2 I26_I24_I2_I0_I0 ( I26_nCv_0n_4_, I26_I24_I2_I0_int_0n[0], I26_I24_I2_I0_int_0n[1] );
  AN2 I26_I25_I2_I0_I2 ( I26_I25_I2_I0_int_0n[0], I26_I25_start, I26_I25_I2_nsel_0n );
  AN2 I26_I25_I2_I0_I1 ( I26_I25_I2_I0_int_0n[1], I26_I25_cv, I26_I25_ha );
  NR2 I26_I25_I2_I0_I0 ( I26_nCv_0n_5_, I26_I25_I2_I0_int_0n[0], I26_I25_I2_I0_int_0n[1] );
  AN2 I26_I26_I2_I0_I2 ( I26_I26_I2_I0_int_0n[0], I26_I26_start, I26_I26_I2_nsel_0n );
  AN2 I26_I26_I2_I0_I1 ( I26_I26_I2_I0_int_0n[1], I26_I26_cv, I26_I26_ha );
  NR2 I26_I26_I2_I0_I0 ( I26_nCv_0n_6_, I26_I26_I2_I0_int_0n[0], I26_I26_I2_I0_int_0n[1] );
  AN2 I26_I27_I2_I0_I2 ( I26_I27_I2_I0_int_0n[0], I26_I27_start, I26_I27_I2_nsel_0n );
  AN2 I26_I27_I2_I0_I1 ( I26_I27_I2_I0_int_0n[1], I26_I27_cv, I26_I27_ha );
  NR2 I26_I27_I2_I0_I0 ( I26_nCv_0n_7_, I26_I27_I2_I0_int_0n[0], I26_I27_I2_I0_int_0n[1] );
  AN2 I26_I28_I2_I0_I2 ( I26_I28_I2_I0_int_0n[0], I26_I28_start, I26_I28_I2_nsel_0n );
  AN2 I26_I28_I2_I0_I1 ( I26_I28_I2_I0_int_0n[1], I26_I28_cv, I26_I28_ha );
  NR2 I26_I28_I2_I0_I0 ( I26_nCv_0n_8_, I26_I28_I2_I0_int_0n[0], I26_I28_I2_I0_int_0n[1] );
  AN2 I26_I29_I2_I0_I2 ( I26_I29_I2_I0_int_0n[0], I26_I29_start, I26_I29_I2_nsel_0n );
  AN2 I26_I29_I2_I0_I1 ( I26_I29_I2_I0_int_0n[1], I26_I29_cv, I26_I29_ha );
  NR2 I26_I29_I2_I0_I0 ( I26_nCv_0n_9_, I26_I29_I2_I0_int_0n[0], I26_I29_I2_I0_int_0n[1] );
  AN2 I26_I30_I2_I0_I2 ( I26_I30_I2_I0_int_0n[0], I26_I30_start, I26_I30_I2_nsel_0n );
  AN2 I26_I30_I2_I0_I1 ( I26_I30_I2_I0_int_0n[1], I26_I30_cv, I26_I30_ha );
  NR2 I26_I30_I2_I0_I0 ( I26_nCv_0n_10_, I26_I30_I2_I0_int_0n[0], I26_I30_I2_I0_int_0n[1] );
  AN2 I26_I31_I2_I0_I2 ( I26_I31_I2_I0_int_0n[0], I26_I31_start, I26_I31_I2_nsel_0n );
  AN2 I26_I31_I2_I0_I1 ( I26_I31_I2_I0_int_0n[1], I26_I31_cv, I26_I31_ha );
  NR2 I26_I31_I2_I0_I0 ( I26_nCv_0n_11_, I26_I31_I2_I0_int_0n[0], I26_I31_I2_I0_int_0n[1] );
  AN2 I26_I32_I2_I0_I2 ( I26_I32_I2_I0_int_0n[0], I26_I32_start, I26_I32_I2_nsel_0n );
  AN2 I26_I32_I2_I0_I1 ( I26_I32_I2_I0_int_0n[1], I26_I32_cv, I26_I32_ha );
  NR2 I26_I32_I2_I0_I0 ( I26_nCv_0n_12_, I26_I32_I2_I0_int_0n[0], I26_I32_I2_I0_int_0n[1] );
  AN2 I26_I33_I2_I0_I2 ( I26_I33_I2_I0_int_0n[0], I26_I33_start, I26_I33_I2_nsel_0n );
  AN2 I26_I33_I2_I0_I1 ( I26_I33_I2_I0_int_0n[1], I26_I33_cv, I26_I33_ha );
  NR2 I26_I33_I2_I0_I0 ( I26_nCv_0n_13_, I26_I33_I2_I0_int_0n[0], I26_I33_I2_I0_int_0n[1] );
  AN2 I26_I34_I2_I0_I2 ( I26_I34_I2_I0_int_0n[0], I26_I34_start, I26_I34_I2_nsel_0n );
  AN2 I26_I34_I2_I0_I1 ( I26_I34_I2_I0_int_0n[1], I26_I34_cv, I26_I34_ha );
  NR2 I26_I34_I2_I0_I0 ( I26_nCv_0n_14_, I26_I34_I2_I0_int_0n[0], I26_I34_I2_I0_int_0n[1] );
  AN2 I26_I35_I2_I0_I2 ( I26_I35_I2_I0_int_0n[0], I26_I35_start, I26_I35_I2_nsel_0n );
  AN2 I26_I35_I2_I0_I1 ( I26_I35_I2_I0_int_0n[1], I26_I35_cv, I26_I35_ha );
  NR2 I26_I35_I2_I0_I0 ( I26_nCv_0n_15_, I26_I35_I2_I0_int_0n[0], I26_I35_I2_I0_int_0n[1] );
  AN2 I26_I36_I2_I0_I2 ( I26_I36_I2_I0_int_0n[0], I26_I36_start, I26_I36_I2_nsel_0n );
  AN2 I26_I36_I2_I0_I1 ( I26_I36_I2_I0_int_0n[1], I26_I36_cv, I26_I36_ha );
  NR2 I26_I36_I2_I0_I0 ( I26_nCv_0n_16_, I26_I36_I2_I0_int_0n[0], I26_I36_I2_I0_int_0n[1] );
  IV I1_I0_I1 ( I1_I0_nsel_0n, I1_select_0n );
  IV I1_I1_I1 ( I1_I1_nsel_0n, I1_select_0n );
  IV I1_I2_I1 ( I1_I2_nsel_0n, I1_select_0n );
  IV I1_I3_I1 ( I1_I3_nsel_0n, I1_select_0n );
  IV I1_I4_I1 ( I1_I4_nsel_0n, I1_select_0n );
  IV I1_I5_I1 ( I1_I5_nsel_0n, I1_select_0n );
  IV I1_I6_I1 ( I1_I6_nsel_0n, I1_select_0n );
  IV I1_I7_I1 ( I1_I7_nsel_0n, I1_select_0n );
  IV I1_I8_I1 ( I1_I8_nsel_0n, I1_select_0n );
  IV I1_I9_I1 ( I1_I9_nsel_0n, I1_select_0n );
  IV I1_I10_I1 ( I1_I10_nsel_0n, I1_select_0n );
  IV I1_I11_I1 ( I1_I11_nsel_0n, I1_select_0n );
  IV I1_I12_I1 ( I1_I12_nsel_0n, I1_select_0n );
  IV I1_I13_I1 ( I1_I13_nsel_0n, I1_select_0n );
  IV I1_I14_I1 ( I1_I14_nsel_0n, I1_select_0n );
  IV I1_I15_I1 ( I1_I15_nsel_0n, I1_select_0n );
  IV I1_I16_I1 ( I1_I16_nsel_0n, I1_select_0n );
  IV I3_I0_I1 ( I3_I0_nsel_0n, I3_select_0n );
  IV I3_I1_I1 ( I3_I1_nsel_0n, I3_select_0n );
  IV I3_I2_I1 ( I3_I2_nsel_0n, I3_select_0n );
  IV I3_I3_I1 ( I3_I3_nsel_0n, I3_select_0n );
  IV I3_I4_I1 ( I3_I4_nsel_0n, I3_select_0n );
  IV I3_I5_I1 ( I3_I5_nsel_0n, I3_select_0n );
  IV I3_I6_I1 ( I3_I6_nsel_0n, I3_select_0n );
  IV I3_I7_I1 ( I3_I7_nsel_0n, I3_select_0n );
  IV I3_I8_I1 ( I3_I8_nsel_0n, I3_select_0n );
  IV I3_I9_I1 ( I3_I9_nsel_0n, I3_select_0n );
  IV I3_I10_I1 ( I3_I10_nsel_0n, I3_select_0n );
  IV I3_I11_I1 ( I3_I11_nsel_0n, I3_select_0n );
  IV I3_I12_I1 ( I3_I12_nsel_0n, I3_select_0n );
  IV I3_I13_I1 ( I3_I13_nsel_0n, I3_select_0n );
  IV I3_I14_I1 ( I3_I14_nsel_0n, I3_select_0n );
  IV I3_I15_I1 ( I3_I15_nsel_0n, I3_select_0n );
  IV I3_I16_I1 ( I3_I16_nsel_0n, I3_select_0n );
  IV I16_I13_I3_I1 ( I16_I13_I3_nsel_0n, I16_I13_ha );
  IV I16_I14_I3_I1 ( I16_I14_I3_nsel_0n, I16_I14_ha );
  IV I16_I15_I3_I1 ( I16_I15_I3_nsel_0n, I16_I15_ha );
  IV I16_I16_I3_I1 ( I16_I16_I3_nsel_0n, I16_I16_ha );
  IV I16_I17_I3_I1 ( I16_I17_I3_nsel_0n, I16_I17_ha );
  IV I16_I18_I3_I1 ( I16_I18_I3_nsel_0n, I16_I18_ha );
  IV I16_I19_I3_I1 ( I16_I19_I3_nsel_0n, I16_I19_ha );
  IV I16_I20_I3_I1 ( I16_I20_I3_nsel_0n, I16_I20_ha );
  IV I16_I21_I3_I1 ( I16_I21_I3_nsel_0n, I16_I21_ha );
  IV I16_I22_I3_I1 ( I16_I22_I3_nsel_0n, I16_I22_ha );
  IV I16_I23_I3_I1 ( I16_I23_I3_nsel_0n, I16_I23_ha );
  IV I16_I24_I3_I1 ( I16_I24_I3_nsel_0n, I16_I24_ha );
  IV I16_I25_I3_I1 ( I16_I25_I3_nsel_0n, I16_I25_ha );
  IV I16_I26_I3_I1 ( I16_I26_I3_nsel_0n, I16_I26_ha );
  IV I16_I27_I3_I1 ( I16_I27_I3_nsel_0n, I16_I27_ha );
  IV I16_I28_I3_I1 ( I16_I28_I3_nsel_0n, I16_I28_ha );
  IV I21_I21_I3_I1 ( I21_I21_I3_nsel_0n, I21_I21_ha );
  IV I21_I22_I3_I1 ( I21_I22_I3_nsel_0n, I21_I22_ha );
  IV I21_I23_I3_I1 ( I21_I23_I3_nsel_0n, I21_I23_ha );
  IV I21_I24_I3_I1 ( I21_I24_I3_nsel_0n, I21_I24_ha );
  IV I21_I25_I3_I1 ( I21_I25_I3_nsel_0n, I21_I25_ha );
  IV I21_I26_I3_I1 ( I21_I26_I3_nsel_0n, I21_I26_ha );
  IV I21_I27_I3_I1 ( I21_I27_I3_nsel_0n, I21_I27_ha );
  IV I21_I28_I3_I1 ( I21_I28_I3_nsel_0n, I21_I28_ha );
  IV I21_I29_I3_I1 ( I21_I29_I3_nsel_0n, I21_I29_ha );
  IV I21_I30_I3_I1 ( I21_I30_I3_nsel_0n, I21_I30_ha );
  IV I21_I31_I3_I1 ( I21_I31_I3_nsel_0n, I21_I31_ha );
  IV I21_I32_I3_I1 ( I21_I32_I3_nsel_0n, I21_I32_ha );
  IV I21_I33_I3_I1 ( I21_I33_I3_nsel_0n, I21_I33_ha );
  IV I21_I34_I3_I1 ( I21_I34_I3_nsel_0n, I21_I34_ha );
  IV I21_I35_I3_I1 ( I21_I35_I3_nsel_0n, I21_I35_ha );
  IV I21_I36_I3_I1 ( I21_I36_I3_nsel_0n, I21_I36_ha );
  IV I26_I21_I3_I1 ( I26_I21_I3_nsel_0n, I26_I21_ha );
  IV I26_I22_I3_I1 ( I26_I22_I3_nsel_0n, I26_I22_ha );
  IV I26_I23_I3_I1 ( I26_I23_I3_nsel_0n, I26_I23_ha );
  IV I26_I24_I3_I1 ( I26_I24_I3_nsel_0n, I26_I24_ha );
  IV I26_I25_I3_I1 ( I26_I25_I3_nsel_0n, I26_I25_ha );
  IV I26_I26_I3_I1 ( I26_I26_I3_nsel_0n, I26_I26_ha );
  IV I26_I27_I3_I1 ( I26_I27_I3_nsel_0n, I26_I27_ha );
  IV I26_I28_I3_I1 ( I26_I28_I3_nsel_0n, I26_I28_ha );
  IV I26_I29_I3_I1 ( I26_I29_I3_nsel_0n, I26_I29_ha );
  IV I26_I30_I3_I1 ( I26_I30_I3_nsel_0n, I26_I30_ha );
  IV I26_I31_I3_I1 ( I26_I31_I3_nsel_0n, I26_I31_ha );
  IV I26_I32_I3_I1 ( I26_I32_I3_nsel_0n, I26_I32_ha );
  IV I26_I33_I3_I1 ( I26_I33_I3_nsel_0n, I26_I33_ha );
  IV I26_I34_I3_I1 ( I26_I34_I3_nsel_0n, I26_I34_ha );
  IV I26_I35_I3_I1 ( I26_I35_I3_nsel_0n, I26_I35_ha );
  IV I26_I36_I3_I1 ( I26_I36_I3_nsel_0n, I26_I36_ha );
  AN2 I1_I0_I0_I2 ( I1_I0_I0_int_0n[0], c24_d[0], I1_I0_nsel_0n );
  AN2 I1_I0_I0_I1 ( I1_I0_I0_int_0n[1], x_0d[0], I1_select_0n );
  OR2 I1_I0_I0_I0 ( c45_d[0], I1_I0_I0_int_0n[0], I1_I0_I0_int_0n[1] );
  AN2 I1_I1_I0_I2 ( I1_I1_I0_int_0n[0], c24_d[1], I1_I1_nsel_0n );
  AN2 I1_I1_I0_I1 ( I1_I1_I0_int_0n[1], x_0d[1], I1_select_0n );
  OR2 I1_I1_I0_I0 ( c45_d[1], I1_I1_I0_int_0n[0], I1_I1_I0_int_0n[1] );
  AN2 I1_I2_I0_I2 ( I1_I2_I0_int_0n[0], c24_d[2], I1_I2_nsel_0n );
  AN2 I1_I2_I0_I1 ( I1_I2_I0_int_0n[1], x_0d[2], I1_select_0n );
  OR2 I1_I2_I0_I0 ( c45_d[2], I1_I2_I0_int_0n[0], I1_I2_I0_int_0n[1] );
  AN2 I1_I3_I0_I2 ( I1_I3_I0_int_0n[0], c24_d[3], I1_I3_nsel_0n );
  AN2 I1_I3_I0_I1 ( I1_I3_I0_int_0n[1], x_0d[3], I1_select_0n );
  OR2 I1_I3_I0_I0 ( c45_d[3], I1_I3_I0_int_0n[0], I1_I3_I0_int_0n[1] );
  AN2 I1_I4_I0_I2 ( I1_I4_I0_int_0n[0], c24_d[4], I1_I4_nsel_0n );
  AN2 I1_I4_I0_I1 ( I1_I4_I0_int_0n[1], x_0d[4], I1_select_0n );
  OR2 I1_I4_I0_I0 ( c45_d[4], I1_I4_I0_int_0n[0], I1_I4_I0_int_0n[1] );
  AN2 I1_I5_I0_I2 ( I1_I5_I0_int_0n[0], c24_d[5], I1_I5_nsel_0n );
  AN2 I1_I5_I0_I1 ( I1_I5_I0_int_0n[1], x_0d[5], I1_select_0n );
  OR2 I1_I5_I0_I0 ( c45_d[5], I1_I5_I0_int_0n[0], I1_I5_I0_int_0n[1] );
  AN2 I1_I6_I0_I2 ( I1_I6_I0_int_0n[0], c24_d[6], I1_I6_nsel_0n );
  AN2 I1_I6_I0_I1 ( I1_I6_I0_int_0n[1], x_0d[6], I1_select_0n );
  OR2 I1_I6_I0_I0 ( c45_d[6], I1_I6_I0_int_0n[0], I1_I6_I0_int_0n[1] );
  AN2 I1_I7_I0_I2 ( I1_I7_I0_int_0n[0], c24_d[7], I1_I7_nsel_0n );
  AN2 I1_I7_I0_I1 ( I1_I7_I0_int_0n[1], x_0d[7], I1_select_0n );
  OR2 I1_I7_I0_I0 ( c45_d[7], I1_I7_I0_int_0n[0], I1_I7_I0_int_0n[1] );
  AN2 I1_I8_I0_I2 ( I1_I8_I0_int_0n[0], c24_d[8], I1_I8_nsel_0n );
  AN2 I1_I8_I0_I1 ( I1_I8_I0_int_0n[1], x_0d[8], I1_select_0n );
  OR2 I1_I8_I0_I0 ( c45_d[8], I1_I8_I0_int_0n[0], I1_I8_I0_int_0n[1] );
  AN2 I1_I9_I0_I2 ( I1_I9_I0_int_0n[0], c24_d[9], I1_I9_nsel_0n );
  AN2 I1_I9_I0_I1 ( I1_I9_I0_int_0n[1], x_0d[9], I1_select_0n );
  OR2 I1_I9_I0_I0 ( c45_d[9], I1_I9_I0_int_0n[0], I1_I9_I0_int_0n[1] );
  AN2 I1_I10_I0_I2 ( I1_I10_I0_int_0n[0], c24_d[10], I1_I10_nsel_0n );
  AN2 I1_I10_I0_I1 ( I1_I10_I0_int_0n[1], x_0d[10], I1_select_0n );
  OR2 I1_I10_I0_I0 ( c45_d[10], I1_I10_I0_int_0n[0], I1_I10_I0_int_0n[1] );
  AN2 I1_I11_I0_I2 ( I1_I11_I0_int_0n[0], c24_d[11], I1_I11_nsel_0n );
  AN2 I1_I11_I0_I1 ( I1_I11_I0_int_0n[1], x_0d[11], I1_select_0n );
  OR2 I1_I11_I0_I0 ( c45_d[11], I1_I11_I0_int_0n[0], I1_I11_I0_int_0n[1] );
  AN2 I1_I12_I0_I2 ( I1_I12_I0_int_0n[0], c24_d[12], I1_I12_nsel_0n );
  AN2 I1_I12_I0_I1 ( I1_I12_I0_int_0n[1], x_0d[12], I1_select_0n );
  OR2 I1_I12_I0_I0 ( c45_d[12], I1_I12_I0_int_0n[0], I1_I12_I0_int_0n[1] );
  AN2 I1_I13_I0_I2 ( I1_I13_I0_int_0n[0], c24_d[13], I1_I13_nsel_0n );
  AN2 I1_I13_I0_I1 ( I1_I13_I0_int_0n[1], x_0d[13], I1_select_0n );
  OR2 I1_I13_I0_I0 ( c45_d[13], I1_I13_I0_int_0n[0], I1_I13_I0_int_0n[1] );
  AN2 I1_I14_I0_I2 ( I1_I14_I0_int_0n[0], c24_d[14], I1_I14_nsel_0n );
  AN2 I1_I14_I0_I1 ( I1_I14_I0_int_0n[1], x_0d[14], I1_select_0n );
  OR2 I1_I14_I0_I0 ( c45_d[14], I1_I14_I0_int_0n[0], I1_I14_I0_int_0n[1] );
  AN2 I1_I15_I0_I2 ( I1_I15_I0_int_0n[0], c24_d[15], I1_I15_nsel_0n );
  AN2 I1_I15_I0_I1 ( I1_I15_I0_int_0n[1], x_0d[15], I1_select_0n );
  OR2 I1_I15_I0_I0 ( c45_d[15], I1_I15_I0_int_0n[0], I1_I15_I0_int_0n[1] );
  AN2 I1_I16_I0_I2 ( I1_I16_I0_int_0n[0], c22_r, I1_I16_nsel_0n );
  AN2 I1_I16_I0_I1 ( I1_I16_I0_int_0n[1], x_0a, I1_select_0n );
  OR2 I1_I16_I0_I0 ( c45_r, I1_I16_I0_int_0n[0], I1_I16_I0_int_0n[1] );
  AN2 I3_I0_I0_I2 ( I3_I0_I0_int_0n[0], c15_d[0], I3_I0_nsel_0n );
  AN2 I3_I0_I0_I1 ( I3_I0_I0_int_0n[1], y_0d[0], I3_select_0n );
  OR2 I3_I0_I0_I0 ( c44_d[0], I3_I0_I0_int_0n[0], I3_I0_I0_int_0n[1] );
  AN2 I3_I1_I0_I2 ( I3_I1_I0_int_0n[0], c15_d[1], I3_I1_nsel_0n );
  AN2 I3_I1_I0_I1 ( I3_I1_I0_int_0n[1], y_0d[1], I3_select_0n );
  OR2 I3_I1_I0_I0 ( c44_d[1], I3_I1_I0_int_0n[0], I3_I1_I0_int_0n[1] );
  AN2 I3_I2_I0_I2 ( I3_I2_I0_int_0n[0], c15_d[2], I3_I2_nsel_0n );
  AN2 I3_I2_I0_I1 ( I3_I2_I0_int_0n[1], y_0d[2], I3_select_0n );
  OR2 I3_I2_I0_I0 ( c44_d[2], I3_I2_I0_int_0n[0], I3_I2_I0_int_0n[1] );
  AN2 I3_I3_I0_I2 ( I3_I3_I0_int_0n[0], c15_d[3], I3_I3_nsel_0n );
  AN2 I3_I3_I0_I1 ( I3_I3_I0_int_0n[1], y_0d[3], I3_select_0n );
  OR2 I3_I3_I0_I0 ( c44_d[3], I3_I3_I0_int_0n[0], I3_I3_I0_int_0n[1] );
  AN2 I3_I4_I0_I2 ( I3_I4_I0_int_0n[0], c15_d[4], I3_I4_nsel_0n );
  AN2 I3_I4_I0_I1 ( I3_I4_I0_int_0n[1], y_0d[4], I3_select_0n );
  OR2 I3_I4_I0_I0 ( c44_d[4], I3_I4_I0_int_0n[0], I3_I4_I0_int_0n[1] );
  AN2 I3_I5_I0_I2 ( I3_I5_I0_int_0n[0], c15_d[5], I3_I5_nsel_0n );
  AN2 I3_I5_I0_I1 ( I3_I5_I0_int_0n[1], y_0d[5], I3_select_0n );
  OR2 I3_I5_I0_I0 ( c44_d[5], I3_I5_I0_int_0n[0], I3_I5_I0_int_0n[1] );
  AN2 I3_I6_I0_I2 ( I3_I6_I0_int_0n[0], c15_d[6], I3_I6_nsel_0n );
  AN2 I3_I6_I0_I1 ( I3_I6_I0_int_0n[1], y_0d[6], I3_select_0n );
  OR2 I3_I6_I0_I0 ( c44_d[6], I3_I6_I0_int_0n[0], I3_I6_I0_int_0n[1] );
  AN2 I3_I7_I0_I2 ( I3_I7_I0_int_0n[0], c15_d[7], I3_I7_nsel_0n );
  AN2 I3_I7_I0_I1 ( I3_I7_I0_int_0n[1], y_0d[7], I3_select_0n );
  OR2 I3_I7_I0_I0 ( c44_d[7], I3_I7_I0_int_0n[0], I3_I7_I0_int_0n[1] );
  AN2 I3_I8_I0_I2 ( I3_I8_I0_int_0n[0], c15_d[8], I3_I8_nsel_0n );
  AN2 I3_I8_I0_I1 ( I3_I8_I0_int_0n[1], y_0d[8], I3_select_0n );
  OR2 I3_I8_I0_I0 ( c44_d[8], I3_I8_I0_int_0n[0], I3_I8_I0_int_0n[1] );
  AN2 I3_I9_I0_I2 ( I3_I9_I0_int_0n[0], c15_d[9], I3_I9_nsel_0n );
  AN2 I3_I9_I0_I1 ( I3_I9_I0_int_0n[1], y_0d[9], I3_select_0n );
  OR2 I3_I9_I0_I0 ( c44_d[9], I3_I9_I0_int_0n[0], I3_I9_I0_int_0n[1] );
  AN2 I3_I10_I0_I2 ( I3_I10_I0_int_0n[0], c15_d[10], I3_I10_nsel_0n );
  AN2 I3_I10_I0_I1 ( I3_I10_I0_int_0n[1], y_0d[10], I3_select_0n );
  OR2 I3_I10_I0_I0 ( c44_d[10], I3_I10_I0_int_0n[0], I3_I10_I0_int_0n[1] );
  AN2 I3_I11_I0_I2 ( I3_I11_I0_int_0n[0], c15_d[11], I3_I11_nsel_0n );
  AN2 I3_I11_I0_I1 ( I3_I11_I0_int_0n[1], y_0d[11], I3_select_0n );
  OR2 I3_I11_I0_I0 ( c44_d[11], I3_I11_I0_int_0n[0], I3_I11_I0_int_0n[1] );
  AN2 I3_I12_I0_I2 ( I3_I12_I0_int_0n[0], c15_d[12], I3_I12_nsel_0n );
  AN2 I3_I12_I0_I1 ( I3_I12_I0_int_0n[1], y_0d[12], I3_select_0n );
  OR2 I3_I12_I0_I0 ( c44_d[12], I3_I12_I0_int_0n[0], I3_I12_I0_int_0n[1] );
  AN2 I3_I13_I0_I2 ( I3_I13_I0_int_0n[0], c15_d[13], I3_I13_nsel_0n );
  AN2 I3_I13_I0_I1 ( I3_I13_I0_int_0n[1], y_0d[13], I3_select_0n );
  OR2 I3_I13_I0_I0 ( c44_d[13], I3_I13_I0_int_0n[0], I3_I13_I0_int_0n[1] );
  AN2 I3_I14_I0_I2 ( I3_I14_I0_int_0n[0], c15_d[14], I3_I14_nsel_0n );
  AN2 I3_I14_I0_I1 ( I3_I14_I0_int_0n[1], y_0d[14], I3_select_0n );
  OR2 I3_I14_I0_I0 ( c44_d[14], I3_I14_I0_int_0n[0], I3_I14_I0_int_0n[1] );
  AN2 I3_I15_I0_I2 ( I3_I15_I0_int_0n[0], c15_d[15], I3_I15_nsel_0n );
  AN2 I3_I15_I0_I1 ( I3_I15_I0_int_0n[1], y_0d[15], I3_select_0n );
  OR2 I3_I15_I0_I0 ( c44_d[15], I3_I15_I0_int_0n[0], I3_I15_I0_int_0n[1] );
  AN2 I3_I16_I0_I2 ( I3_I16_I0_int_0n[0], c13_r, I3_I16_nsel_0n );
  AN2 I3_I16_I0_I1 ( I3_I16_I0_int_0n[1], y_0a, I3_select_0n );
  OR2 I3_I16_I0_I0 ( c44_r, I3_I16_I0_int_0n[0], I3_I16_I0_int_0n[1] );
  AN2 I16_I13_I3_I0_I2 ( I16_I13_I3_I0_int_0n[0], I16_n_0n[0], I16_I13_I3_nsel_0n );
  AN2 I16_I13_I3_I0_I1 ( I16_I13_I3_I0_int_0n[1], I16_vcc, I16_I13_ha );
  OR2 I16_I13_I3_I0_I0 ( I16_c_0n_1_, I16_I13_I3_I0_int_0n[0], I16_I13_I3_I0_int_0n[1] );
  AN2 I16_I14_I3_I0_I2 ( I16_I14_I3_I0_int_0n[0], I16_n_0n[1], I16_I14_I3_nsel_0n );
  AN2 I16_I14_I3_I0_I1 ( I16_I14_I3_I0_int_0n[1], I16_c_0n_1_, I16_I14_ha );
  OR2 I16_I14_I3_I0_I0 ( I16_c_0n_2_, I16_I14_I3_I0_int_0n[0], I16_I14_I3_I0_int_0n[1] );
  AN2 I16_I15_I3_I0_I2 ( I16_I15_I3_I0_int_0n[0], I16_n_0n[2], I16_I15_I3_nsel_0n );
  AN2 I16_I15_I3_I0_I1 ( I16_I15_I3_I0_int_0n[1], I16_c_0n_2_, I16_I15_ha );
  OR2 I16_I15_I3_I0_I0 ( I16_c_0n_3_, I16_I15_I3_I0_int_0n[0], I16_I15_I3_I0_int_0n[1] );
  AN2 I16_I16_I3_I0_I2 ( I16_I16_I3_I0_int_0n[0], I16_n_0n[3], I16_I16_I3_nsel_0n );
  AN2 I16_I16_I3_I0_I1 ( I16_I16_I3_I0_int_0n[1], I16_c_0n_3_, I16_I16_ha );
  OR2 I16_I16_I3_I0_I0 ( I16_c_0n_4_, I16_I16_I3_I0_int_0n[0], I16_I16_I3_I0_int_0n[1] );
  AN2 I16_I17_I3_I0_I2 ( I16_I17_I3_I0_int_0n[0], I16_n_0n[4], I16_I17_I3_nsel_0n );
  AN2 I16_I17_I3_I0_I1 ( I16_I17_I3_I0_int_0n[1], I16_c_0n_4_, I16_I17_ha );
  OR2 I16_I17_I3_I0_I0 ( I16_c_0n_5_, I16_I17_I3_I0_int_0n[0], I16_I17_I3_I0_int_0n[1] );
  AN2 I16_I18_I3_I0_I2 ( I16_I18_I3_I0_int_0n[0], I16_n_0n[5], I16_I18_I3_nsel_0n );
  AN2 I16_I18_I3_I0_I1 ( I16_I18_I3_I0_int_0n[1], I16_c_0n_5_, I16_I18_ha );
  OR2 I16_I18_I3_I0_I0 ( I16_c_0n_6_, I16_I18_I3_I0_int_0n[0], I16_I18_I3_I0_int_0n[1] );
  AN2 I16_I19_I3_I0_I2 ( I16_I19_I3_I0_int_0n[0], I16_n_0n[6], I16_I19_I3_nsel_0n );
  AN2 I16_I19_I3_I0_I1 ( I16_I19_I3_I0_int_0n[1], I16_c_0n_6_, I16_I19_ha );
  OR2 I16_I19_I3_I0_I0 ( I16_c_0n_7_, I16_I19_I3_I0_int_0n[0], I16_I19_I3_I0_int_0n[1] );
  AN2 I16_I20_I3_I0_I2 ( I16_I20_I3_I0_int_0n[0], I16_n_0n[7], I16_I20_I3_nsel_0n );
  AN2 I16_I20_I3_I0_I1 ( I16_I20_I3_I0_int_0n[1], I16_c_0n_7_, I16_I20_ha );
  OR2 I16_I20_I3_I0_I0 ( I16_c_0n_8_, I16_I20_I3_I0_int_0n[0], I16_I20_I3_I0_int_0n[1] );
  AN2 I16_I21_I3_I0_I2 ( I16_I21_I3_I0_int_0n[0], I16_n_0n[8], I16_I21_I3_nsel_0n );
  AN2 I16_I21_I3_I0_I1 ( I16_I21_I3_I0_int_0n[1], I16_c_0n_8_, I16_I21_ha );
  OR2 I16_I21_I3_I0_I0 ( I16_c_0n_9_, I16_I21_I3_I0_int_0n[0], I16_I21_I3_I0_int_0n[1] );
  AN2 I16_I22_I3_I0_I2 ( I16_I22_I3_I0_int_0n[0], I16_n_0n[9], I16_I22_I3_nsel_0n );
  AN2 I16_I22_I3_I0_I1 ( I16_I22_I3_I0_int_0n[1], I16_c_0n_9_, I16_I22_ha );
  OR2 I16_I22_I3_I0_I0 ( I16_c_0n_10_, I16_I22_I3_I0_int_0n[0], I16_I22_I3_I0_int_0n[1] );
  AN2 I16_I23_I3_I0_I2 ( I16_I23_I3_I0_int_0n[0], I16_n_0n[10], I16_I23_I3_nsel_0n );
  AN2 I16_I23_I3_I0_I1 ( I16_I23_I3_I0_int_0n[1], I16_c_0n_10_, I16_I23_ha );
  OR2 I16_I23_I3_I0_I0 ( I16_c_0n_11_, I16_I23_I3_I0_int_0n[0], I16_I23_I3_I0_int_0n[1] );
  AN2 I16_I24_I3_I0_I2 ( I16_I24_I3_I0_int_0n[0], I16_n_0n[11], I16_I24_I3_nsel_0n );
  AN2 I16_I24_I3_I0_I1 ( I16_I24_I3_I0_int_0n[1], I16_c_0n_11_, I16_I24_ha );
  OR2 I16_I24_I3_I0_I0 ( I16_c_0n_12_, I16_I24_I3_I0_int_0n[0], I16_I24_I3_I0_int_0n[1] );
  AN2 I16_I25_I3_I0_I2 ( I16_I25_I3_I0_int_0n[0], I16_n_0n[12], I16_I25_I3_nsel_0n );
  AN2 I16_I25_I3_I0_I1 ( I16_I25_I3_I0_int_0n[1], I16_c_0n_12_, I16_I25_ha );
  OR2 I16_I25_I3_I0_I0 ( I16_c_0n_13_, I16_I25_I3_I0_int_0n[0], I16_I25_I3_I0_int_0n[1] );
  AN2 I16_I26_I3_I0_I2 ( I16_I26_I3_I0_int_0n[0], I16_n_0n[13], I16_I26_I3_nsel_0n );
  AN2 I16_I26_I3_I0_I1 ( I16_I26_I3_I0_int_0n[1], I16_c_0n_13_, I16_I26_ha );
  OR2 I16_I26_I3_I0_I0 ( I16_c_0n_14_, I16_I26_I3_I0_int_0n[0], I16_I26_I3_I0_int_0n[1] );
  AN2 I16_I27_I3_I0_I2 ( I16_I27_I3_I0_int_0n[0], I16_n_0n[14], I16_I27_I3_nsel_0n );
  AN2 I16_I27_I3_I0_I1 ( I16_I27_I3_I0_int_0n[1], I16_c_0n_14_, I16_I27_ha );
  OR2 I16_I27_I3_I0_I0 ( I16_c_0n_15_, I16_I27_I3_I0_int_0n[0], I16_I27_I3_I0_int_0n[1] );
  AN2 I16_I28_I3_I0_I2 ( I16_I28_I3_I0_int_0n[0], I16_n_0n[15], I16_I28_I3_nsel_0n );
  AN2 I16_I28_I3_I0_I1 ( I16_I28_I3_I0_int_0n[1], I16_c_0n_15_, I16_I28_ha );
  OR2 I16_I28_I3_I0_I0 ( I16_c_0n_16_, I16_I28_I3_I0_int_0n[0], I16_I28_I3_I0_int_0n[1] );
  AN2 I21_I21_I3_I0_I2 ( I21_I21_I3_I0_int_0n[0], I21_n_0n[0], I21_I21_I3_nsel_0n );
  AN2 I21_I21_I3_I0_I1 ( I21_I21_I3_I0_int_0n[1], I21_vcc, I21_I21_ha );
  OR2 I21_I21_I3_I0_I0 ( I21_c_0n[1], I21_I21_I3_I0_int_0n[0], I21_I21_I3_I0_int_0n[1] );
  AN2 I21_I22_I3_I0_I2 ( I21_I22_I3_I0_int_0n[0], I21_n_0n[1], I21_I22_I3_nsel_0n );
  AN2 I21_I22_I3_I0_I1 ( I21_I22_I3_I0_int_0n[1], I21_c_0n[1], I21_I22_ha );
  OR2 I21_I22_I3_I0_I0 ( I21_c_0n[2], I21_I22_I3_I0_int_0n[0], I21_I22_I3_I0_int_0n[1] );
  AN2 I21_I23_I3_I0_I2 ( I21_I23_I3_I0_int_0n[0], I21_n_0n[2], I21_I23_I3_nsel_0n );
  AN2 I21_I23_I3_I0_I1 ( I21_I23_I3_I0_int_0n[1], I21_c_0n[2], I21_I23_ha );
  OR2 I21_I23_I3_I0_I0 ( I21_c_0n[3], I21_I23_I3_I0_int_0n[0], I21_I23_I3_I0_int_0n[1] );
  AN2 I21_I24_I3_I0_I2 ( I21_I24_I3_I0_int_0n[0], I21_n_0n[3], I21_I24_I3_nsel_0n );
  AN2 I21_I24_I3_I0_I1 ( I21_I24_I3_I0_int_0n[1], I21_c_0n[3], I21_I24_ha );
  OR2 I21_I24_I3_I0_I0 ( I21_c_0n[4], I21_I24_I3_I0_int_0n[0], I21_I24_I3_I0_int_0n[1] );
  AN2 I21_I25_I3_I0_I2 ( I21_I25_I3_I0_int_0n[0], I21_n_0n[4], I21_I25_I3_nsel_0n );
  AN2 I21_I25_I3_I0_I1 ( I21_I25_I3_I0_int_0n[1], I21_c_0n[4], I21_I25_ha );
  OR2 I21_I25_I3_I0_I0 ( I21_c_0n[5], I21_I25_I3_I0_int_0n[0], I21_I25_I3_I0_int_0n[1] );
  AN2 I21_I26_I3_I0_I2 ( I21_I26_I3_I0_int_0n[0], I21_n_0n[5], I21_I26_I3_nsel_0n );
  AN2 I21_I26_I3_I0_I1 ( I21_I26_I3_I0_int_0n[1], I21_c_0n[5], I21_I26_ha );
  OR2 I21_I26_I3_I0_I0 ( I21_c_0n[6], I21_I26_I3_I0_int_0n[0], I21_I26_I3_I0_int_0n[1] );
  AN2 I21_I27_I3_I0_I2 ( I21_I27_I3_I0_int_0n[0], I21_n_0n[6], I21_I27_I3_nsel_0n );
  AN2 I21_I27_I3_I0_I1 ( I21_I27_I3_I0_int_0n[1], I21_c_0n[6], I21_I27_ha );
  OR2 I21_I27_I3_I0_I0 ( I21_c_0n[7], I21_I27_I3_I0_int_0n[0], I21_I27_I3_I0_int_0n[1] );
  AN2 I21_I28_I3_I0_I2 ( I21_I28_I3_I0_int_0n[0], I21_n_0n[7], I21_I28_I3_nsel_0n );
  AN2 I21_I28_I3_I0_I1 ( I21_I28_I3_I0_int_0n[1], I21_c_0n[7], I21_I28_ha );
  OR2 I21_I28_I3_I0_I0 ( I21_c_0n[8], I21_I28_I3_I0_int_0n[0], I21_I28_I3_I0_int_0n[1] );
  AN2 I21_I29_I3_I0_I2 ( I21_I29_I3_I0_int_0n[0], I21_n_0n[8], I21_I29_I3_nsel_0n );
  AN2 I21_I29_I3_I0_I1 ( I21_I29_I3_I0_int_0n[1], I21_c_0n[8], I21_I29_ha );
  OR2 I21_I29_I3_I0_I0 ( I21_c_0n[9], I21_I29_I3_I0_int_0n[0], I21_I29_I3_I0_int_0n[1] );
  AN2 I21_I30_I3_I0_I2 ( I21_I30_I3_I0_int_0n[0], I21_n_0n[9], I21_I30_I3_nsel_0n );
  AN2 I21_I30_I3_I0_I1 ( I21_I30_I3_I0_int_0n[1], I21_c_0n[9], I21_I30_ha );
  OR2 I21_I30_I3_I0_I0 ( I21_c_0n[10], I21_I30_I3_I0_int_0n[0], I21_I30_I3_I0_int_0n[1] );
  AN2 I21_I31_I3_I0_I2 ( I21_I31_I3_I0_int_0n[0], I21_n_0n[10], I21_I31_I3_nsel_0n );
  AN2 I21_I31_I3_I0_I1 ( I21_I31_I3_I0_int_0n[1], I21_c_0n[10], I21_I31_ha );
  OR2 I21_I31_I3_I0_I0 ( I21_c_0n[11], I21_I31_I3_I0_int_0n[0], I21_I31_I3_I0_int_0n[1] );
  AN2 I21_I32_I3_I0_I2 ( I21_I32_I3_I0_int_0n[0], I21_n_0n[11], I21_I32_I3_nsel_0n );
  AN2 I21_I32_I3_I0_I1 ( I21_I32_I3_I0_int_0n[1], I21_c_0n[11], I21_I32_ha );
  OR2 I21_I32_I3_I0_I0 ( I21_c_0n[12], I21_I32_I3_I0_int_0n[0], I21_I32_I3_I0_int_0n[1] );
  AN2 I21_I33_I3_I0_I2 ( I21_I33_I3_I0_int_0n[0], I21_n_0n[12], I21_I33_I3_nsel_0n );
  AN2 I21_I33_I3_I0_I1 ( I21_I33_I3_I0_int_0n[1], I21_c_0n[12], I21_I33_ha );
  OR2 I21_I33_I3_I0_I0 ( I21_c_0n[13], I21_I33_I3_I0_int_0n[0], I21_I33_I3_I0_int_0n[1] );
  AN2 I21_I34_I3_I0_I2 ( I21_I34_I3_I0_int_0n[0], I21_n_0n[13], I21_I34_I3_nsel_0n );
  AN2 I21_I34_I3_I0_I1 ( I21_I34_I3_I0_int_0n[1], I21_c_0n[13], I21_I34_ha );
  OR2 I21_I34_I3_I0_I0 ( I21_c_0n[14], I21_I34_I3_I0_int_0n[0], I21_I34_I3_I0_int_0n[1] );
  AN2 I21_I35_I3_I0_I2 ( I21_I35_I3_I0_int_0n[0], I21_n_0n[14], I21_I35_I3_nsel_0n );
  AN2 I21_I35_I3_I0_I1 ( I21_I35_I3_I0_int_0n[1], I21_c_0n[14], I21_I35_ha );
  OR2 I21_I35_I3_I0_I0 ( I21_c_0n[15], I21_I35_I3_I0_int_0n[0], I21_I35_I3_I0_int_0n[1] );
  AN2 I21_I36_I3_I0_I2 ( I21_I36_I3_I0_int_0n[0], I21_n_0n[15], I21_I36_I3_nsel_0n );
  AN2 I21_I36_I3_I0_I1 ( I21_I36_I3_I0_int_0n[1], I21_c_0n[15], I21_I36_ha );
  OR2 I21_I36_I3_I0_I0 ( I21_c_0n[16], I21_I36_I3_I0_int_0n[0], I21_I36_I3_I0_int_0n[1] );
  AN2 I26_I21_I3_I0_I2 ( I26_I21_I3_I0_int_0n[0], I26_n_0n[0], I26_I21_I3_nsel_0n );
  AN2 I26_I21_I3_I0_I1 ( I26_I21_I3_I0_int_0n[1], I26_vcc, I26_I21_ha );
  OR2 I26_I21_I3_I0_I0 ( I26_c_0n[1], I26_I21_I3_I0_int_0n[0], I26_I21_I3_I0_int_0n[1] );
  AN2 I26_I22_I3_I0_I2 ( I26_I22_I3_I0_int_0n[0], I26_n_0n[1], I26_I22_I3_nsel_0n );
  AN2 I26_I22_I3_I0_I1 ( I26_I22_I3_I0_int_0n[1], I26_c_0n[1], I26_I22_ha );
  OR2 I26_I22_I3_I0_I0 ( I26_c_0n[2], I26_I22_I3_I0_int_0n[0], I26_I22_I3_I0_int_0n[1] );
  AN2 I26_I23_I3_I0_I2 ( I26_I23_I3_I0_int_0n[0], I26_n_0n[2], I26_I23_I3_nsel_0n );
  AN2 I26_I23_I3_I0_I1 ( I26_I23_I3_I0_int_0n[1], I26_c_0n[2], I26_I23_ha );
  OR2 I26_I23_I3_I0_I0 ( I26_c_0n[3], I26_I23_I3_I0_int_0n[0], I26_I23_I3_I0_int_0n[1] );
  AN2 I26_I24_I3_I0_I2 ( I26_I24_I3_I0_int_0n[0], I26_n_0n[3], I26_I24_I3_nsel_0n );
  AN2 I26_I24_I3_I0_I1 ( I26_I24_I3_I0_int_0n[1], I26_c_0n[3], I26_I24_ha );
  OR2 I26_I24_I3_I0_I0 ( I26_c_0n[4], I26_I24_I3_I0_int_0n[0], I26_I24_I3_I0_int_0n[1] );
  AN2 I26_I25_I3_I0_I2 ( I26_I25_I3_I0_int_0n[0], I26_n_0n[4], I26_I25_I3_nsel_0n );
  AN2 I26_I25_I3_I0_I1 ( I26_I25_I3_I0_int_0n[1], I26_c_0n[4], I26_I25_ha );
  OR2 I26_I25_I3_I0_I0 ( I26_c_0n[5], I26_I25_I3_I0_int_0n[0], I26_I25_I3_I0_int_0n[1] );
  AN2 I26_I26_I3_I0_I2 ( I26_I26_I3_I0_int_0n[0], I26_n_0n[5], I26_I26_I3_nsel_0n );
  AN2 I26_I26_I3_I0_I1 ( I26_I26_I3_I0_int_0n[1], I26_c_0n[5], I26_I26_ha );
  OR2 I26_I26_I3_I0_I0 ( I26_c_0n[6], I26_I26_I3_I0_int_0n[0], I26_I26_I3_I0_int_0n[1] );
  AN2 I26_I27_I3_I0_I2 ( I26_I27_I3_I0_int_0n[0], I26_n_0n[6], I26_I27_I3_nsel_0n );
  AN2 I26_I27_I3_I0_I1 ( I26_I27_I3_I0_int_0n[1], I26_c_0n[6], I26_I27_ha );
  OR2 I26_I27_I3_I0_I0 ( I26_c_0n[7], I26_I27_I3_I0_int_0n[0], I26_I27_I3_I0_int_0n[1] );
  AN2 I26_I28_I3_I0_I2 ( I26_I28_I3_I0_int_0n[0], I26_n_0n[7], I26_I28_I3_nsel_0n );
  AN2 I26_I28_I3_I0_I1 ( I26_I28_I3_I0_int_0n[1], I26_c_0n[7], I26_I28_ha );
  OR2 I26_I28_I3_I0_I0 ( I26_c_0n[8], I26_I28_I3_I0_int_0n[0], I26_I28_I3_I0_int_0n[1] );
  AN2 I26_I29_I3_I0_I2 ( I26_I29_I3_I0_int_0n[0], I26_n_0n[8], I26_I29_I3_nsel_0n );
  AN2 I26_I29_I3_I0_I1 ( I26_I29_I3_I0_int_0n[1], I26_c_0n[8], I26_I29_ha );
  OR2 I26_I29_I3_I0_I0 ( I26_c_0n[9], I26_I29_I3_I0_int_0n[0], I26_I29_I3_I0_int_0n[1] );
  AN2 I26_I30_I3_I0_I2 ( I26_I30_I3_I0_int_0n[0], I26_n_0n[9], I26_I30_I3_nsel_0n );
  AN2 I26_I30_I3_I0_I1 ( I26_I30_I3_I0_int_0n[1], I26_c_0n[9], I26_I30_ha );
  OR2 I26_I30_I3_I0_I0 ( I26_c_0n[10], I26_I30_I3_I0_int_0n[0], I26_I30_I3_I0_int_0n[1] );
  AN2 I26_I31_I3_I0_I2 ( I26_I31_I3_I0_int_0n[0], I26_n_0n[10], I26_I31_I3_nsel_0n );
  AN2 I26_I31_I3_I0_I1 ( I26_I31_I3_I0_int_0n[1], I26_c_0n[10], I26_I31_ha );
  OR2 I26_I31_I3_I0_I0 ( I26_c_0n[11], I26_I31_I3_I0_int_0n[0], I26_I31_I3_I0_int_0n[1] );
  AN2 I26_I32_I3_I0_I2 ( I26_I32_I3_I0_int_0n[0], I26_n_0n[11], I26_I32_I3_nsel_0n );
  AN2 I26_I32_I3_I0_I1 ( I26_I32_I3_I0_int_0n[1], I26_c_0n[11], I26_I32_ha );
  OR2 I26_I32_I3_I0_I0 ( I26_c_0n[12], I26_I32_I3_I0_int_0n[0], I26_I32_I3_I0_int_0n[1] );
  AN2 I26_I33_I3_I0_I2 ( I26_I33_I3_I0_int_0n[0], I26_n_0n[12], I26_I33_I3_nsel_0n );
  AN2 I26_I33_I3_I0_I1 ( I26_I33_I3_I0_int_0n[1], I26_c_0n[12], I26_I33_ha );
  OR2 I26_I33_I3_I0_I0 ( I26_c_0n[13], I26_I33_I3_I0_int_0n[0], I26_I33_I3_I0_int_0n[1] );
  AN2 I26_I34_I3_I0_I2 ( I26_I34_I3_I0_int_0n[0], I26_n_0n[13], I26_I34_I3_nsel_0n );
  AN2 I26_I34_I3_I0_I1 ( I26_I34_I3_I0_int_0n[1], I26_c_0n[13], I26_I34_ha );
  OR2 I26_I34_I3_I0_I0 ( I26_c_0n[14], I26_I34_I3_I0_int_0n[0], I26_I34_I3_I0_int_0n[1] );
  AN2 I26_I35_I3_I0_I2 ( I26_I35_I3_I0_int_0n[0], I26_n_0n[14], I26_I35_I3_nsel_0n );
  AN2 I26_I35_I3_I0_I1 ( I26_I35_I3_I0_int_0n[1], I26_c_0n[14], I26_I35_ha );
  OR2 I26_I35_I3_I0_I0 ( I26_c_0n[15], I26_I35_I3_I0_int_0n[0], I26_I35_I3_I0_int_0n[1] );
  AN2 I26_I36_I3_I0_I2 ( I26_I36_I3_I0_int_0n[0], I26_n_0n[15], I26_I36_I3_nsel_0n );
  AN2 I26_I36_I3_I0_I1 ( I26_I36_I3_I0_int_0n[1], I26_c_0n[15], I26_I36_ha );
  OR2 I26_I36_I3_I0_I0 ( I26_c_0n[16], I26_I36_I3_I0_int_0n[0], I26_I36_I3_I0_int_0n[1] );
endmodule

/*
    `booth_mul16.v'
    Balsa Verilog netlist file
    Created: Tue Jan 14 14:23:22 JST 2014
    By: xaos@kikurage (Linux)
    With net-verilog (balsa-netlist) version: 4.0
    Using technology: aclass/four_b_rb
    Command line : (balsa-netlist -Xaclass booth_mul16)

    Using `propagate-globals'
    The design contains no global nets
*/

module buf1 (
  z,
  a
);
  output z;
  input a;
  wire na_0n;
  IV I0 (z, na_0n);
  IV I1 (na_0n, a);
endmodule

module BrzAdapt_33_17_s5_false_s5_false (
  out_0r, out_0a, out_0d,
  inp_0r, inp_0a, inp_0d
);
  input out_0r;
  output out_0a;
  output [32:0] out_0d;
  output inp_0r;
  input inp_0a;
  input [16:0] inp_0d;
  wire extend_0n;
  wire gnd;
  GND gnd_cell_instance (gnd);
  assign out_0a = inp_0a;
  assign inp_0r = out_0r;
  assign out_0d[17] = gnd;
  assign out_0d[18] = gnd;
  assign out_0d[19] = gnd;
  assign out_0d[20] = gnd;
  assign out_0d[21] = gnd;
  assign out_0d[22] = gnd;
  assign out_0d[23] = gnd;
  assign out_0d[24] = gnd;
  assign out_0d[25] = gnd;
  assign out_0d[26] = gnd;
  assign out_0d[27] = gnd;
  assign out_0d[28] = gnd;
  assign out_0d[29] = gnd;
  assign out_0d[30] = gnd;
  assign out_0d[31] = gnd;
  assign out_0d[32] = gnd;
  assign out_0d[0] = inp_0d[0];
  assign out_0d[1] = inp_0d[1];
  assign out_0d[2] = inp_0d[2];
  assign out_0d[3] = inp_0d[3];
  assign out_0d[4] = inp_0d[4];
  assign out_0d[5] = inp_0d[5];
  assign out_0d[6] = inp_0d[6];
  assign out_0d[7] = inp_0d[7];
  assign out_0d[8] = inp_0d[8];
  assign out_0d[9] = inp_0d[9];
  assign out_0d[10] = inp_0d[10];
  assign out_0d[11] = inp_0d[11];
  assign out_0d[12] = inp_0d[12];
  assign out_0d[13] = inp_0d[13];
  assign out_0d[14] = inp_0d[14];
  assign out_0d[15] = inp_0d[15];
  assign out_0d[16] = inp_0d[16];
endmodule

module demux2 (
  i,
  o0,
  o1,
  s
);
  input i;
  output o0;
  output o1;
  input s;
  wire ns_0n;
  AN2 I0 (o1, i, s);
  AN2 I1 (o0, i, ns_0n);
  IV I2 (ns_0n, s);
endmodule

module BrzBar_2 (
  guard_0r, guard_0a, guard_0d,
  activate_0r, activate_0a,
  guardInput_0r, guardInput_0a, guardInput_0d,
  guardInput_1r, guardInput_1a, guardInput_1d,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a
);
  input guard_0r;
  output guard_0a;
  output guard_0d;
  input activate_0r;
  output activate_0a;
  output guardInput_0r;
  input guardInput_0a;
  input guardInput_0d;
  output guardInput_1r;
  input guardInput_1a;
  input guardInput_1d;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  wire [2:0] bypass_0n;
  wire [1:0] outReq_0n;
  C2 I0 (activateOut_0r, activate_0r, outReq_0n[0]);
  C2 I1 (activateOut_1r, activate_0r, outReq_0n[1]);
  demux2 I2 (bypass_0n[0], bypass_0n[1], outReq_0n[0], guardInput_0d);
  demux2 I3 (bypass_0n[1], bypass_0n[2], outReq_0n[1], guardInput_1d);
  assign bypass_0n[0] = activate_0r;
  OR3 I5 (activate_0a, activateOut_0a, activateOut_1a, bypass_0n[2]);
  OR2 I6 (guard_0d, guardInput_0d, guardInput_1d);
  C2 I7 (guard_0a, guardInput_0a, guardInput_1a);
  assign guardInput_0r = guard_0r;
  assign guardInput_1r = guard_0r;
endmodule

module BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m (
  out_0r, out_0a, out_0d,
  inpA_0r, inpA_0a, inpA_0d,
  inpB_0r, inpB_0a, inpB_0d
);
  input out_0r;
  output out_0a;
  output out_0d;
  output inpA_0r;
  input inpA_0a;
  input inpA_0d;
  output inpB_0r;
  input inpB_0a;
  input inpB_0d;
  wire start_0n;
  wire nStart_0n;
  wire [1:0] nCv_0n;
  wire [1:0] c_0n;
  wire eq_0n;
  wire addOut_0n;
  wire w_0n;
  wire n_0n;
  wire v_0n;
  wire z_0n;
  wire nz_0n;
  wire nxv_0n;
  wire done_0n;
  AN2 I0 (out_0d, n_0n, w_0n);
  assign done_0n = start_0n;
  assign n_0n = inpB_0d;
  assign w_0n = inpA_0d;
  assign out_0a = done_0n;
  C2 I5 (start_0n, inpA_0a, inpB_0a);
  assign inpA_0r = out_0r;
  assign inpB_0r = out_0r;
endmodule

module ao22 (
  q,
  i0,
  i1,
  i2,
  i3
);
  output q;
  input i0;
  input i1;
  input i2;
  input i3;
  wire [1:0] int_0n;
  OR2 I0 (q, int_0n[0], int_0n[1]);
  AN2 I1 (int_0n[1], i2, i3);
  AN2 I2 (int_0n[0], i0, i1);
endmodule

module mux2 (
  out,
  in0,
  in1,
  sel
);
  output out;
  input in0;
  input in1;
  input sel;
  wire nsel_0n;
  ao22 I0 (out, in0, nsel_0n, in1, sel);
  IV I1 (nsel_0n, sel);
endmodule

module aoi22 (
  q,
  i0,
  i1,
  i2,
  i3
);
  output q;
  input i0;
  input i1;
  input i2;
  input i3;
  wire [1:0] int_0n;
  NR2 I0 (q, int_0n[0], int_0n[1]);
  AN2 I1 (int_0n[1], i2, i3);
  AN2 I2 (int_0n[0], i0, i1);
endmodule

module nmux2 (
  out,
  in0,
  in1,
  sel
);
  output out;
  input in0;
  input in1;
  input sel;
  wire nsel_0n;
  aoi22 I0 (out, in0, nsel_0n, in1, sel);
  IV I1 (nsel_0n, sel);
endmodule

module balsa_fa (
  nStart,
  A,
  B,
  nCVi,
  Ci,
  nCVo,
  Co,
  sum
);
  input nStart;
  input A;
  input B;
  input nCVi;
  input Ci;
  output nCVo;
  output Co;
  output sum;
  wire start;
  wire ha;
  wire cv;
  IV I0 (start, nStart);
  NR2 I1 (cv, nStart, nCVi);
  nmux2 I2 (nCVo, start, cv, ha);
  mux2 I3 (Co, A, Ci, ha);
  EO I4 (ha, A, B);
  EO I5 (sum, ha, Ci);
endmodule

module BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m (
  out_0r, out_0a, out_0d,
  inpA_0r, inpA_0a, inpA_0d,
  inpB_0r, inpB_0a, inpB_0d
);
  input out_0r;
  output out_0a;
  output [33:0] out_0d;
  output inpA_0r;
  input inpA_0a;
  input [32:0] inpA_0d;
  output inpB_0r;
  input inpB_0a;
  input [32:0] inpB_0d;
  wire [11:0] internal_0n;
  wire start_0n;
  wire nStart_0n;
  wire [33:0] nCv_0n;
  wire [33:0] c_0n;
  wire [32:0] eq_0n;
  wire [32:0] addOut_0n;
  wire [32:0] w_0n;
  wire [32:0] n_0n;
  wire v_0n;
  wire z_0n;
  wire nz_0n;
  wire nxv_0n;
  wire done_0n;
  wire gnd;
  GND gnd_cell_instance (gnd);
  NR4 I0 (internal_0n[0], nCv_0n[1], nCv_0n[2], nCv_0n[3], nCv_0n[4]);
  NR4 I1 (internal_0n[1], nCv_0n[5], nCv_0n[6], nCv_0n[7], nCv_0n[8]);
  NR4 I2 (internal_0n[2], nCv_0n[9], nCv_0n[10], nCv_0n[11], nCv_0n[12]);
  NR4 I3 (internal_0n[3], nCv_0n[13], nCv_0n[14], nCv_0n[15], nCv_0n[16]);
  NR4 I4 (internal_0n[4], nCv_0n[17], nCv_0n[18], nCv_0n[19], nCv_0n[20]);
  NR4 I5 (internal_0n[5], nCv_0n[21], nCv_0n[22], nCv_0n[23], nCv_0n[24]);
  NR4 I6 (internal_0n[6], nCv_0n[25], nCv_0n[26], nCv_0n[27], nCv_0n[28]);
  NR2 I7 (internal_0n[7], nCv_0n[29], nCv_0n[30]);
  NR3 I8 (internal_0n[8], nCv_0n[31], nCv_0n[32], nCv_0n[33]);
  ND4 I9 (internal_0n[9], internal_0n[0], internal_0n[1], internal_0n[2], internal_0n[3]);
  ND2 I10 (internal_0n[10], internal_0n[4], internal_0n[5]);
  ND3 I11 (internal_0n[11], internal_0n[6], internal_0n[7], internal_0n[8]);
  NR3 I12 (done_0n, internal_0n[9], internal_0n[10], internal_0n[11]);
  assign out_0d[0] = addOut_0n[0];
  assign out_0d[1] = addOut_0n[1];
  assign out_0d[2] = addOut_0n[2];
  assign out_0d[3] = addOut_0n[3];
  assign out_0d[4] = addOut_0n[4];
  assign out_0d[5] = addOut_0n[5];
  assign out_0d[6] = addOut_0n[6];
  assign out_0d[7] = addOut_0n[7];
  assign out_0d[8] = addOut_0n[8];
  assign out_0d[9] = addOut_0n[9];
  assign out_0d[10] = addOut_0n[10];
  assign out_0d[11] = addOut_0n[11];
  assign out_0d[12] = addOut_0n[12];
  assign out_0d[13] = addOut_0n[13];
  assign out_0d[14] = addOut_0n[14];
  assign out_0d[15] = addOut_0n[15];
  assign out_0d[16] = addOut_0n[16];
  assign out_0d[17] = addOut_0n[17];
  assign out_0d[18] = addOut_0n[18];
  assign out_0d[19] = addOut_0n[19];
  assign out_0d[20] = addOut_0n[20];
  assign out_0d[21] = addOut_0n[21];
  assign out_0d[22] = addOut_0n[22];
  assign out_0d[23] = addOut_0n[23];
  assign out_0d[24] = addOut_0n[24];
  assign out_0d[25] = addOut_0n[25];
  assign out_0d[26] = addOut_0n[26];
  assign out_0d[27] = addOut_0n[27];
  assign out_0d[28] = addOut_0n[28];
  assign out_0d[29] = addOut_0n[29];
  assign out_0d[30] = addOut_0n[30];
  assign out_0d[31] = addOut_0n[31];
  assign out_0d[32] = addOut_0n[32];
  assign out_0d[33] = c_0n[33];
  balsa_fa I47 (nStart_0n, n_0n[0], w_0n[0], nCv_0n[0], c_0n[0], nCv_0n[1], c_0n[1], addOut_0n[0]);
  balsa_fa I48 (nStart_0n, n_0n[1], w_0n[1], nCv_0n[1], c_0n[1], nCv_0n[2], c_0n[2], addOut_0n[1]);
  balsa_fa I49 (nStart_0n, n_0n[2], w_0n[2], nCv_0n[2], c_0n[2], nCv_0n[3], c_0n[3], addOut_0n[2]);
  balsa_fa I50 (nStart_0n, n_0n[3], w_0n[3], nCv_0n[3], c_0n[3], nCv_0n[4], c_0n[4], addOut_0n[3]);
  balsa_fa I51 (nStart_0n, n_0n[4], w_0n[4], nCv_0n[4], c_0n[4], nCv_0n[5], c_0n[5], addOut_0n[4]);
  balsa_fa I52 (nStart_0n, n_0n[5], w_0n[5], nCv_0n[5], c_0n[5], nCv_0n[6], c_0n[6], addOut_0n[5]);
  balsa_fa I53 (nStart_0n, n_0n[6], w_0n[6], nCv_0n[6], c_0n[6], nCv_0n[7], c_0n[7], addOut_0n[6]);
  balsa_fa I54 (nStart_0n, n_0n[7], w_0n[7], nCv_0n[7], c_0n[7], nCv_0n[8], c_0n[8], addOut_0n[7]);
  balsa_fa I55 (nStart_0n, n_0n[8], w_0n[8], nCv_0n[8], c_0n[8], nCv_0n[9], c_0n[9], addOut_0n[8]);
  balsa_fa I56 (nStart_0n, n_0n[9], w_0n[9], nCv_0n[9], c_0n[9], nCv_0n[10], c_0n[10], addOut_0n[9]);
  balsa_fa I57 (nStart_0n, n_0n[10], w_0n[10], nCv_0n[10], c_0n[10], nCv_0n[11], c_0n[11], addOut_0n[10]);
  balsa_fa I58 (nStart_0n, n_0n[11], w_0n[11], nCv_0n[11], c_0n[11], nCv_0n[12], c_0n[12], addOut_0n[11]);
  balsa_fa I59 (nStart_0n, n_0n[12], w_0n[12], nCv_0n[12], c_0n[12], nCv_0n[13], c_0n[13], addOut_0n[12]);
  balsa_fa I60 (nStart_0n, n_0n[13], w_0n[13], nCv_0n[13], c_0n[13], nCv_0n[14], c_0n[14], addOut_0n[13]);
  balsa_fa I61 (nStart_0n, n_0n[14], w_0n[14], nCv_0n[14], c_0n[14], nCv_0n[15], c_0n[15], addOut_0n[14]);
  balsa_fa I62 (nStart_0n, n_0n[15], w_0n[15], nCv_0n[15], c_0n[15], nCv_0n[16], c_0n[16], addOut_0n[15]);
  balsa_fa I63 (nStart_0n, n_0n[16], w_0n[16], nCv_0n[16], c_0n[16], nCv_0n[17], c_0n[17], addOut_0n[16]);
  balsa_fa I64 (nStart_0n, n_0n[17], w_0n[17], nCv_0n[17], c_0n[17], nCv_0n[18], c_0n[18], addOut_0n[17]);
  balsa_fa I65 (nStart_0n, n_0n[18], w_0n[18], nCv_0n[18], c_0n[18], nCv_0n[19], c_0n[19], addOut_0n[18]);
  balsa_fa I66 (nStart_0n, n_0n[19], w_0n[19], nCv_0n[19], c_0n[19], nCv_0n[20], c_0n[20], addOut_0n[19]);
  balsa_fa I67 (nStart_0n, n_0n[20], w_0n[20], nCv_0n[20], c_0n[20], nCv_0n[21], c_0n[21], addOut_0n[20]);
  balsa_fa I68 (nStart_0n, n_0n[21], w_0n[21], nCv_0n[21], c_0n[21], nCv_0n[22], c_0n[22], addOut_0n[21]);
  balsa_fa I69 (nStart_0n, n_0n[22], w_0n[22], nCv_0n[22], c_0n[22], nCv_0n[23], c_0n[23], addOut_0n[22]);
  balsa_fa I70 (nStart_0n, n_0n[23], w_0n[23], nCv_0n[23], c_0n[23], nCv_0n[24], c_0n[24], addOut_0n[23]);
  balsa_fa I71 (nStart_0n, n_0n[24], w_0n[24], nCv_0n[24], c_0n[24], nCv_0n[25], c_0n[25], addOut_0n[24]);
  balsa_fa I72 (nStart_0n, n_0n[25], w_0n[25], nCv_0n[25], c_0n[25], nCv_0n[26], c_0n[26], addOut_0n[25]);
  balsa_fa I73 (nStart_0n, n_0n[26], w_0n[26], nCv_0n[26], c_0n[26], nCv_0n[27], c_0n[27], addOut_0n[26]);
  balsa_fa I74 (nStart_0n, n_0n[27], w_0n[27], nCv_0n[27], c_0n[27], nCv_0n[28], c_0n[28], addOut_0n[27]);
  balsa_fa I75 (nStart_0n, n_0n[28], w_0n[28], nCv_0n[28], c_0n[28], nCv_0n[29], c_0n[29], addOut_0n[28]);
  balsa_fa I76 (nStart_0n, n_0n[29], w_0n[29], nCv_0n[29], c_0n[29], nCv_0n[30], c_0n[30], addOut_0n[29]);
  balsa_fa I77 (nStart_0n, n_0n[30], w_0n[30], nCv_0n[30], c_0n[30], nCv_0n[31], c_0n[31], addOut_0n[30]);
  balsa_fa I78 (nStart_0n, n_0n[31], w_0n[31], nCv_0n[31], c_0n[31], nCv_0n[32], c_0n[32], addOut_0n[31]);
  balsa_fa I79 (nStart_0n, n_0n[32], w_0n[32], nCv_0n[32], c_0n[32], nCv_0n[33], c_0n[33], addOut_0n[32]);
  assign nCv_0n[0] = nStart_0n;
  assign c_0n[0] = gnd;
  IV I82 (nStart_0n, start_0n);
  assign n_0n[0] = inpB_0d[0];
  assign n_0n[1] = inpB_0d[1];
  assign n_0n[2] = inpB_0d[2];
  assign n_0n[3] = inpB_0d[3];
  assign n_0n[4] = inpB_0d[4];
  assign n_0n[5] = inpB_0d[5];
  assign n_0n[6] = inpB_0d[6];
  assign n_0n[7] = inpB_0d[7];
  assign n_0n[8] = inpB_0d[8];
  assign n_0n[9] = inpB_0d[9];
  assign n_0n[10] = inpB_0d[10];
  assign n_0n[11] = inpB_0d[11];
  assign n_0n[12] = inpB_0d[12];
  assign n_0n[13] = inpB_0d[13];
  assign n_0n[14] = inpB_0d[14];
  assign n_0n[15] = inpB_0d[15];
  assign n_0n[16] = inpB_0d[16];
  assign n_0n[17] = inpB_0d[17];
  assign n_0n[18] = inpB_0d[18];
  assign n_0n[19] = inpB_0d[19];
  assign n_0n[20] = inpB_0d[20];
  assign n_0n[21] = inpB_0d[21];
  assign n_0n[22] = inpB_0d[22];
  assign n_0n[23] = inpB_0d[23];
  assign n_0n[24] = inpB_0d[24];
  assign n_0n[25] = inpB_0d[25];
  assign n_0n[26] = inpB_0d[26];
  assign n_0n[27] = inpB_0d[27];
  assign n_0n[28] = inpB_0d[28];
  assign n_0n[29] = inpB_0d[29];
  assign n_0n[30] = inpB_0d[30];
  assign n_0n[31] = inpB_0d[31];
  assign n_0n[32] = inpB_0d[32];
  assign w_0n[0] = inpA_0d[0];
  assign w_0n[1] = inpA_0d[1];
  assign w_0n[2] = inpA_0d[2];
  assign w_0n[3] = inpA_0d[3];
  assign w_0n[4] = inpA_0d[4];
  assign w_0n[5] = inpA_0d[5];
  assign w_0n[6] = inpA_0d[6];
  assign w_0n[7] = inpA_0d[7];
  assign w_0n[8] = inpA_0d[8];
  assign w_0n[9] = inpA_0d[9];
  assign w_0n[10] = inpA_0d[10];
  assign w_0n[11] = inpA_0d[11];
  assign w_0n[12] = inpA_0d[12];
  assign w_0n[13] = inpA_0d[13];
  assign w_0n[14] = inpA_0d[14];
  assign w_0n[15] = inpA_0d[15];
  assign w_0n[16] = inpA_0d[16];
  assign w_0n[17] = inpA_0d[17];
  assign w_0n[18] = inpA_0d[18];
  assign w_0n[19] = inpA_0d[19];
  assign w_0n[20] = inpA_0d[20];
  assign w_0n[21] = inpA_0d[21];
  assign w_0n[22] = inpA_0d[22];
  assign w_0n[23] = inpA_0d[23];
  assign w_0n[24] = inpA_0d[24];
  assign w_0n[25] = inpA_0d[25];
  assign w_0n[26] = inpA_0d[26];
  assign w_0n[27] = inpA_0d[27];
  assign w_0n[28] = inpA_0d[28];
  assign w_0n[29] = inpA_0d[29];
  assign w_0n[30] = inpA_0d[30];
  assign w_0n[31] = inpA_0d[31];
  assign w_0n[32] = inpA_0d[32];
  assign out_0a = done_0n;
  C2 I150 (start_0n, inpA_0a, inpB_0a);
  assign inpA_0r = out_0r;
  assign inpB_0r = out_0r;
endmodule

module BrzCallMux_33_49 (
  inp_0r, inp_0a, inp_0d,
  inp_1r, inp_1a, inp_1d,
  inp_2r, inp_2a, inp_2d,
  inp_3r, inp_3a, inp_3d,
  inp_4r, inp_4a, inp_4d,
  inp_5r, inp_5a, inp_5d,
  inp_6r, inp_6a, inp_6d,
  inp_7r, inp_7a, inp_7d,
  inp_8r, inp_8a, inp_8d,
  inp_9r, inp_9a, inp_9d,
  inp_10r, inp_10a, inp_10d,
  inp_11r, inp_11a, inp_11d,
  inp_12r, inp_12a, inp_12d,
  inp_13r, inp_13a, inp_13d,
  inp_14r, inp_14a, inp_14d,
  inp_15r, inp_15a, inp_15d,
  inp_16r, inp_16a, inp_16d,
  inp_17r, inp_17a, inp_17d,
  inp_18r, inp_18a, inp_18d,
  inp_19r, inp_19a, inp_19d,
  inp_20r, inp_20a, inp_20d,
  inp_21r, inp_21a, inp_21d,
  inp_22r, inp_22a, inp_22d,
  inp_23r, inp_23a, inp_23d,
  inp_24r, inp_24a, inp_24d,
  inp_25r, inp_25a, inp_25d,
  inp_26r, inp_26a, inp_26d,
  inp_27r, inp_27a, inp_27d,
  inp_28r, inp_28a, inp_28d,
  inp_29r, inp_29a, inp_29d,
  inp_30r, inp_30a, inp_30d,
  inp_31r, inp_31a, inp_31d,
  inp_32r, inp_32a, inp_32d,
  inp_33r, inp_33a, inp_33d,
  inp_34r, inp_34a, inp_34d,
  inp_35r, inp_35a, inp_35d,
  inp_36r, inp_36a, inp_36d,
  inp_37r, inp_37a, inp_37d,
  inp_38r, inp_38a, inp_38d,
  inp_39r, inp_39a, inp_39d,
  inp_40r, inp_40a, inp_40d,
  inp_41r, inp_41a, inp_41d,
  inp_42r, inp_42a, inp_42d,
  inp_43r, inp_43a, inp_43d,
  inp_44r, inp_44a, inp_44d,
  inp_45r, inp_45a, inp_45d,
  inp_46r, inp_46a, inp_46d,
  inp_47r, inp_47a, inp_47d,
  inp_48r, inp_48a, inp_48d,
  out_0r, out_0a, out_0d
);
  input inp_0r;
  output inp_0a;
  input [32:0] inp_0d;
  input inp_1r;
  output inp_1a;
  input [32:0] inp_1d;
  input inp_2r;
  output inp_2a;
  input [32:0] inp_2d;
  input inp_3r;
  output inp_3a;
  input [32:0] inp_3d;
  input inp_4r;
  output inp_4a;
  input [32:0] inp_4d;
  input inp_5r;
  output inp_5a;
  input [32:0] inp_5d;
  input inp_6r;
  output inp_6a;
  input [32:0] inp_6d;
  input inp_7r;
  output inp_7a;
  input [32:0] inp_7d;
  input inp_8r;
  output inp_8a;
  input [32:0] inp_8d;
  input inp_9r;
  output inp_9a;
  input [32:0] inp_9d;
  input inp_10r;
  output inp_10a;
  input [32:0] inp_10d;
  input inp_11r;
  output inp_11a;
  input [32:0] inp_11d;
  input inp_12r;
  output inp_12a;
  input [32:0] inp_12d;
  input inp_13r;
  output inp_13a;
  input [32:0] inp_13d;
  input inp_14r;
  output inp_14a;
  input [32:0] inp_14d;
  input inp_15r;
  output inp_15a;
  input [32:0] inp_15d;
  input inp_16r;
  output inp_16a;
  input [32:0] inp_16d;
  input inp_17r;
  output inp_17a;
  input [32:0] inp_17d;
  input inp_18r;
  output inp_18a;
  input [32:0] inp_18d;
  input inp_19r;
  output inp_19a;
  input [32:0] inp_19d;
  input inp_20r;
  output inp_20a;
  input [32:0] inp_20d;
  input inp_21r;
  output inp_21a;
  input [32:0] inp_21d;
  input inp_22r;
  output inp_22a;
  input [32:0] inp_22d;
  input inp_23r;
  output inp_23a;
  input [32:0] inp_23d;
  input inp_24r;
  output inp_24a;
  input [32:0] inp_24d;
  input inp_25r;
  output inp_25a;
  input [32:0] inp_25d;
  input inp_26r;
  output inp_26a;
  input [32:0] inp_26d;
  input inp_27r;
  output inp_27a;
  input [32:0] inp_27d;
  input inp_28r;
  output inp_28a;
  input [32:0] inp_28d;
  input inp_29r;
  output inp_29a;
  input [32:0] inp_29d;
  input inp_30r;
  output inp_30a;
  input [32:0] inp_30d;
  input inp_31r;
  output inp_31a;
  input [32:0] inp_31d;
  input inp_32r;
  output inp_32a;
  input [32:0] inp_32d;
  input inp_33r;
  output inp_33a;
  input [32:0] inp_33d;
  input inp_34r;
  output inp_34a;
  input [32:0] inp_34d;
  input inp_35r;
  output inp_35a;
  input [32:0] inp_35d;
  input inp_36r;
  output inp_36a;
  input [32:0] inp_36d;
  input inp_37r;
  output inp_37a;
  input [32:0] inp_37d;
  input inp_38r;
  output inp_38a;
  input [32:0] inp_38d;
  input inp_39r;
  output inp_39a;
  input [32:0] inp_39d;
  input inp_40r;
  output inp_40a;
  input [32:0] inp_40d;
  input inp_41r;
  output inp_41a;
  input [32:0] inp_41d;
  input inp_42r;
  output inp_42a;
  input [32:0] inp_42d;
  input inp_43r;
  output inp_43a;
  input [32:0] inp_43d;
  input inp_44r;
  output inp_44a;
  input [32:0] inp_44d;
  input inp_45r;
  output inp_45a;
  input [32:0] inp_45d;
  input inp_46r;
  output inp_46a;
  input [32:0] inp_46d;
  input inp_47r;
  output inp_47a;
  input [32:0] inp_47d;
  input inp_48r;
  output inp_48a;
  input [32:0] inp_48d;
  output out_0r;
  input out_0a;
  output [32:0] out_0d;
  wire [577:0] internal_0n;
  wire [32:0] muxOut_0n;
  wire select_0n;
  wire nselect_0n;
  wire [48:0] nwaySelect_0n;
  wire [32:0] nwayMuxOut_0n;
  wire [32:0] nwayMuxOut_1n;
  wire [32:0] nwayMuxOut_2n;
  wire [32:0] nwayMuxOut_3n;
  wire [32:0] nwayMuxOut_4n;
  wire [32:0] nwayMuxOut_5n;
  wire [32:0] nwayMuxOut_6n;
  wire [32:0] nwayMuxOut_7n;
  wire [32:0] nwayMuxOut_8n;
  wire [32:0] nwayMuxOut_9n;
  wire [32:0] nwayMuxOut_10n;
  wire [32:0] nwayMuxOut_11n;
  wire [32:0] nwayMuxOut_12n;
  wire [32:0] nwayMuxOut_13n;
  wire [32:0] nwayMuxOut_14n;
  wire [32:0] nwayMuxOut_15n;
  wire [32:0] nwayMuxOut_16n;
  wire [32:0] nwayMuxOut_17n;
  wire [32:0] nwayMuxOut_18n;
  wire [32:0] nwayMuxOut_19n;
  wire [32:0] nwayMuxOut_20n;
  wire [32:0] nwayMuxOut_21n;
  wire [32:0] nwayMuxOut_22n;
  wire [32:0] nwayMuxOut_23n;
  wire [32:0] nwayMuxOut_24n;
  wire [32:0] nwayMuxOut_25n;
  wire [32:0] nwayMuxOut_26n;
  wire [32:0] nwayMuxOut_27n;
  wire [32:0] nwayMuxOut_28n;
  wire [32:0] nwayMuxOut_29n;
  wire [32:0] nwayMuxOut_30n;
  wire [32:0] nwayMuxOut_31n;
  wire [32:0] nwayMuxOut_32n;
  wire [32:0] nwayMuxOut_33n;
  wire [32:0] nwayMuxOut_34n;
  wire [32:0] nwayMuxOut_35n;
  wire [32:0] nwayMuxOut_36n;
  wire [32:0] nwayMuxOut_37n;
  wire [32:0] nwayMuxOut_38n;
  wire [32:0] nwayMuxOut_39n;
  wire [32:0] nwayMuxOut_40n;
  wire [32:0] nwayMuxOut_41n;
  wire [32:0] nwayMuxOut_42n;
  wire [32:0] nwayMuxOut_43n;
  wire [32:0] nwayMuxOut_44n;
  wire [32:0] nwayMuxOut_45n;
  wire [32:0] nwayMuxOut_46n;
  wire [32:0] nwayMuxOut_47n;
  wire [32:0] nwayMuxOut_48n;
  ND4 I0 (internal_0n[0], nwayMuxOut_0n[0], nwayMuxOut_1n[0], nwayMuxOut_2n[0], nwayMuxOut_3n[0]);
  ND4 I1 (internal_0n[1], nwayMuxOut_4n[0], nwayMuxOut_5n[0], nwayMuxOut_6n[0], nwayMuxOut_7n[0]);
  ND4 I2 (internal_0n[2], nwayMuxOut_8n[0], nwayMuxOut_9n[0], nwayMuxOut_10n[0], nwayMuxOut_11n[0]);
  ND4 I3 (internal_0n[3], nwayMuxOut_12n[0], nwayMuxOut_13n[0], nwayMuxOut_14n[0], nwayMuxOut_15n[0]);
  ND4 I4 (internal_0n[4], nwayMuxOut_16n[0], nwayMuxOut_17n[0], nwayMuxOut_18n[0], nwayMuxOut_19n[0]);
  ND4 I5 (internal_0n[5], nwayMuxOut_20n[0], nwayMuxOut_21n[0], nwayMuxOut_22n[0], nwayMuxOut_23n[0]);
  ND4 I6 (internal_0n[6], nwayMuxOut_24n[0], nwayMuxOut_25n[0], nwayMuxOut_26n[0], nwayMuxOut_27n[0]);
  ND4 I7 (internal_0n[7], nwayMuxOut_28n[0], nwayMuxOut_29n[0], nwayMuxOut_30n[0], nwayMuxOut_31n[0]);
  ND4 I8 (internal_0n[8], nwayMuxOut_32n[0], nwayMuxOut_33n[0], nwayMuxOut_34n[0], nwayMuxOut_35n[0]);
  ND4 I9 (internal_0n[9], nwayMuxOut_36n[0], nwayMuxOut_37n[0], nwayMuxOut_38n[0], nwayMuxOut_39n[0]);
  ND4 I10 (internal_0n[10], nwayMuxOut_40n[0], nwayMuxOut_41n[0], nwayMuxOut_42n[0], nwayMuxOut_43n[0]);
  ND2 I11 (internal_0n[11], nwayMuxOut_44n[0], nwayMuxOut_45n[0]);
  ND3 I12 (internal_0n[12], nwayMuxOut_46n[0], nwayMuxOut_47n[0], nwayMuxOut_48n[0]);
  NR4 I13 (internal_0n[13], internal_0n[0], internal_0n[1], internal_0n[2], internal_0n[3]);
  NR4 I14 (internal_0n[14], internal_0n[4], internal_0n[5], internal_0n[6], internal_0n[7]);
  NR2 I15 (internal_0n[15], internal_0n[8], internal_0n[9]);
  NR3 I16 (internal_0n[16], internal_0n[10], internal_0n[11], internal_0n[12]);
  ND4 I17 (out_0d[0], internal_0n[13], internal_0n[14], internal_0n[15], internal_0n[16]);
  ND4 I18 (internal_0n[17], nwayMuxOut_0n[1], nwayMuxOut_1n[1], nwayMuxOut_2n[1], nwayMuxOut_3n[1]);
  ND4 I19 (internal_0n[18], nwayMuxOut_4n[1], nwayMuxOut_5n[1], nwayMuxOut_6n[1], nwayMuxOut_7n[1]);
  ND4 I20 (internal_0n[19], nwayMuxOut_8n[1], nwayMuxOut_9n[1], nwayMuxOut_10n[1], nwayMuxOut_11n[1]);
  ND4 I21 (internal_0n[20], nwayMuxOut_12n[1], nwayMuxOut_13n[1], nwayMuxOut_14n[1], nwayMuxOut_15n[1]);
  ND4 I22 (internal_0n[21], nwayMuxOut_16n[1], nwayMuxOut_17n[1], nwayMuxOut_18n[1], nwayMuxOut_19n[1]);
  ND4 I23 (internal_0n[22], nwayMuxOut_20n[1], nwayMuxOut_21n[1], nwayMuxOut_22n[1], nwayMuxOut_23n[1]);
  ND4 I24 (internal_0n[23], nwayMuxOut_24n[1], nwayMuxOut_25n[1], nwayMuxOut_26n[1], nwayMuxOut_27n[1]);
  ND4 I25 (internal_0n[24], nwayMuxOut_28n[1], nwayMuxOut_29n[1], nwayMuxOut_30n[1], nwayMuxOut_31n[1]);
  ND4 I26 (internal_0n[25], nwayMuxOut_32n[1], nwayMuxOut_33n[1], nwayMuxOut_34n[1], nwayMuxOut_35n[1]);
  ND4 I27 (internal_0n[26], nwayMuxOut_36n[1], nwayMuxOut_37n[1], nwayMuxOut_38n[1], nwayMuxOut_39n[1]);
  ND4 I28 (internal_0n[27], nwayMuxOut_40n[1], nwayMuxOut_41n[1], nwayMuxOut_42n[1], nwayMuxOut_43n[1]);
  ND2 I29 (internal_0n[28], nwayMuxOut_44n[1], nwayMuxOut_45n[1]);
  ND3 I30 (internal_0n[29], nwayMuxOut_46n[1], nwayMuxOut_47n[1], nwayMuxOut_48n[1]);
  NR4 I31 (internal_0n[30], internal_0n[17], internal_0n[18], internal_0n[19], internal_0n[20]);
  NR4 I32 (internal_0n[31], internal_0n[21], internal_0n[22], internal_0n[23], internal_0n[24]);
  NR2 I33 (internal_0n[32], internal_0n[25], internal_0n[26]);
  NR3 I34 (internal_0n[33], internal_0n[27], internal_0n[28], internal_0n[29]);
  ND4 I35 (out_0d[1], internal_0n[30], internal_0n[31], internal_0n[32], internal_0n[33]);
  ND4 I36 (internal_0n[34], nwayMuxOut_0n[2], nwayMuxOut_1n[2], nwayMuxOut_2n[2], nwayMuxOut_3n[2]);
  ND4 I37 (internal_0n[35], nwayMuxOut_4n[2], nwayMuxOut_5n[2], nwayMuxOut_6n[2], nwayMuxOut_7n[2]);
  ND4 I38 (internal_0n[36], nwayMuxOut_8n[2], nwayMuxOut_9n[2], nwayMuxOut_10n[2], nwayMuxOut_11n[2]);
  ND4 I39 (internal_0n[37], nwayMuxOut_12n[2], nwayMuxOut_13n[2], nwayMuxOut_14n[2], nwayMuxOut_15n[2]);
  ND4 I40 (internal_0n[38], nwayMuxOut_16n[2], nwayMuxOut_17n[2], nwayMuxOut_18n[2], nwayMuxOut_19n[2]);
  ND4 I41 (internal_0n[39], nwayMuxOut_20n[2], nwayMuxOut_21n[2], nwayMuxOut_22n[2], nwayMuxOut_23n[2]);
  ND4 I42 (internal_0n[40], nwayMuxOut_24n[2], nwayMuxOut_25n[2], nwayMuxOut_26n[2], nwayMuxOut_27n[2]);
  ND4 I43 (internal_0n[41], nwayMuxOut_28n[2], nwayMuxOut_29n[2], nwayMuxOut_30n[2], nwayMuxOut_31n[2]);
  ND4 I44 (internal_0n[42], nwayMuxOut_32n[2], nwayMuxOut_33n[2], nwayMuxOut_34n[2], nwayMuxOut_35n[2]);
  ND4 I45 (internal_0n[43], nwayMuxOut_36n[2], nwayMuxOut_37n[2], nwayMuxOut_38n[2], nwayMuxOut_39n[2]);
  ND4 I46 (internal_0n[44], nwayMuxOut_40n[2], nwayMuxOut_41n[2], nwayMuxOut_42n[2], nwayMuxOut_43n[2]);
  ND2 I47 (internal_0n[45], nwayMuxOut_44n[2], nwayMuxOut_45n[2]);
  ND3 I48 (internal_0n[46], nwayMuxOut_46n[2], nwayMuxOut_47n[2], nwayMuxOut_48n[2]);
  NR4 I49 (internal_0n[47], internal_0n[34], internal_0n[35], internal_0n[36], internal_0n[37]);
  NR4 I50 (internal_0n[48], internal_0n[38], internal_0n[39], internal_0n[40], internal_0n[41]);
  NR2 I51 (internal_0n[49], internal_0n[42], internal_0n[43]);
  NR3 I52 (internal_0n[50], internal_0n[44], internal_0n[45], internal_0n[46]);
  ND4 I53 (out_0d[2], internal_0n[47], internal_0n[48], internal_0n[49], internal_0n[50]);
  ND4 I54 (internal_0n[51], nwayMuxOut_0n[3], nwayMuxOut_1n[3], nwayMuxOut_2n[3], nwayMuxOut_3n[3]);
  ND4 I55 (internal_0n[52], nwayMuxOut_4n[3], nwayMuxOut_5n[3], nwayMuxOut_6n[3], nwayMuxOut_7n[3]);
  ND4 I56 (internal_0n[53], nwayMuxOut_8n[3], nwayMuxOut_9n[3], nwayMuxOut_10n[3], nwayMuxOut_11n[3]);
  ND4 I57 (internal_0n[54], nwayMuxOut_12n[3], nwayMuxOut_13n[3], nwayMuxOut_14n[3], nwayMuxOut_15n[3]);
  ND4 I58 (internal_0n[55], nwayMuxOut_16n[3], nwayMuxOut_17n[3], nwayMuxOut_18n[3], nwayMuxOut_19n[3]);
  ND4 I59 (internal_0n[56], nwayMuxOut_20n[3], nwayMuxOut_21n[3], nwayMuxOut_22n[3], nwayMuxOut_23n[3]);
  ND4 I60 (internal_0n[57], nwayMuxOut_24n[3], nwayMuxOut_25n[3], nwayMuxOut_26n[3], nwayMuxOut_27n[3]);
  ND4 I61 (internal_0n[58], nwayMuxOut_28n[3], nwayMuxOut_29n[3], nwayMuxOut_30n[3], nwayMuxOut_31n[3]);
  ND4 I62 (internal_0n[59], nwayMuxOut_32n[3], nwayMuxOut_33n[3], nwayMuxOut_34n[3], nwayMuxOut_35n[3]);
  ND4 I63 (internal_0n[60], nwayMuxOut_36n[3], nwayMuxOut_37n[3], nwayMuxOut_38n[3], nwayMuxOut_39n[3]);
  ND4 I64 (internal_0n[61], nwayMuxOut_40n[3], nwayMuxOut_41n[3], nwayMuxOut_42n[3], nwayMuxOut_43n[3]);
  ND2 I65 (internal_0n[62], nwayMuxOut_44n[3], nwayMuxOut_45n[3]);
  ND3 I66 (internal_0n[63], nwayMuxOut_46n[3], nwayMuxOut_47n[3], nwayMuxOut_48n[3]);
  NR4 I67 (internal_0n[64], internal_0n[51], internal_0n[52], internal_0n[53], internal_0n[54]);
  NR4 I68 (internal_0n[65], internal_0n[55], internal_0n[56], internal_0n[57], internal_0n[58]);
  NR2 I69 (internal_0n[66], internal_0n[59], internal_0n[60]);
  NR3 I70 (internal_0n[67], internal_0n[61], internal_0n[62], internal_0n[63]);
  ND4 I71 (out_0d[3], internal_0n[64], internal_0n[65], internal_0n[66], internal_0n[67]);
  ND4 I72 (internal_0n[68], nwayMuxOut_0n[4], nwayMuxOut_1n[4], nwayMuxOut_2n[4], nwayMuxOut_3n[4]);
  ND4 I73 (internal_0n[69], nwayMuxOut_4n[4], nwayMuxOut_5n[4], nwayMuxOut_6n[4], nwayMuxOut_7n[4]);
  ND4 I74 (internal_0n[70], nwayMuxOut_8n[4], nwayMuxOut_9n[4], nwayMuxOut_10n[4], nwayMuxOut_11n[4]);
  ND4 I75 (internal_0n[71], nwayMuxOut_12n[4], nwayMuxOut_13n[4], nwayMuxOut_14n[4], nwayMuxOut_15n[4]);
  ND4 I76 (internal_0n[72], nwayMuxOut_16n[4], nwayMuxOut_17n[4], nwayMuxOut_18n[4], nwayMuxOut_19n[4]);
  ND4 I77 (internal_0n[73], nwayMuxOut_20n[4], nwayMuxOut_21n[4], nwayMuxOut_22n[4], nwayMuxOut_23n[4]);
  ND4 I78 (internal_0n[74], nwayMuxOut_24n[4], nwayMuxOut_25n[4], nwayMuxOut_26n[4], nwayMuxOut_27n[4]);
  ND4 I79 (internal_0n[75], nwayMuxOut_28n[4], nwayMuxOut_29n[4], nwayMuxOut_30n[4], nwayMuxOut_31n[4]);
  ND4 I80 (internal_0n[76], nwayMuxOut_32n[4], nwayMuxOut_33n[4], nwayMuxOut_34n[4], nwayMuxOut_35n[4]);
  ND4 I81 (internal_0n[77], nwayMuxOut_36n[4], nwayMuxOut_37n[4], nwayMuxOut_38n[4], nwayMuxOut_39n[4]);
  ND4 I82 (internal_0n[78], nwayMuxOut_40n[4], nwayMuxOut_41n[4], nwayMuxOut_42n[4], nwayMuxOut_43n[4]);
  ND2 I83 (internal_0n[79], nwayMuxOut_44n[4], nwayMuxOut_45n[4]);
  ND3 I84 (internal_0n[80], nwayMuxOut_46n[4], nwayMuxOut_47n[4], nwayMuxOut_48n[4]);
  NR4 I85 (internal_0n[81], internal_0n[68], internal_0n[69], internal_0n[70], internal_0n[71]);
  NR4 I86 (internal_0n[82], internal_0n[72], internal_0n[73], internal_0n[74], internal_0n[75]);
  NR2 I87 (internal_0n[83], internal_0n[76], internal_0n[77]);
  NR3 I88 (internal_0n[84], internal_0n[78], internal_0n[79], internal_0n[80]);
  ND4 I89 (out_0d[4], internal_0n[81], internal_0n[82], internal_0n[83], internal_0n[84]);
  ND4 I90 (internal_0n[85], nwayMuxOut_0n[5], nwayMuxOut_1n[5], nwayMuxOut_2n[5], nwayMuxOut_3n[5]);
  ND4 I91 (internal_0n[86], nwayMuxOut_4n[5], nwayMuxOut_5n[5], nwayMuxOut_6n[5], nwayMuxOut_7n[5]);
  ND4 I92 (internal_0n[87], nwayMuxOut_8n[5], nwayMuxOut_9n[5], nwayMuxOut_10n[5], nwayMuxOut_11n[5]);
  ND4 I93 (internal_0n[88], nwayMuxOut_12n[5], nwayMuxOut_13n[5], nwayMuxOut_14n[5], nwayMuxOut_15n[5]);
  ND4 I94 (internal_0n[89], nwayMuxOut_16n[5], nwayMuxOut_17n[5], nwayMuxOut_18n[5], nwayMuxOut_19n[5]);
  ND4 I95 (internal_0n[90], nwayMuxOut_20n[5], nwayMuxOut_21n[5], nwayMuxOut_22n[5], nwayMuxOut_23n[5]);
  ND4 I96 (internal_0n[91], nwayMuxOut_24n[5], nwayMuxOut_25n[5], nwayMuxOut_26n[5], nwayMuxOut_27n[5]);
  ND4 I97 (internal_0n[92], nwayMuxOut_28n[5], nwayMuxOut_29n[5], nwayMuxOut_30n[5], nwayMuxOut_31n[5]);
  ND4 I98 (internal_0n[93], nwayMuxOut_32n[5], nwayMuxOut_33n[5], nwayMuxOut_34n[5], nwayMuxOut_35n[5]);
  ND4 I99 (internal_0n[94], nwayMuxOut_36n[5], nwayMuxOut_37n[5], nwayMuxOut_38n[5], nwayMuxOut_39n[5]);
  ND4 I100 (internal_0n[95], nwayMuxOut_40n[5], nwayMuxOut_41n[5], nwayMuxOut_42n[5], nwayMuxOut_43n[5]);
  ND2 I101 (internal_0n[96], nwayMuxOut_44n[5], nwayMuxOut_45n[5]);
  ND3 I102 (internal_0n[97], nwayMuxOut_46n[5], nwayMuxOut_47n[5], nwayMuxOut_48n[5]);
  NR4 I103 (internal_0n[98], internal_0n[85], internal_0n[86], internal_0n[87], internal_0n[88]);
  NR4 I104 (internal_0n[99], internal_0n[89], internal_0n[90], internal_0n[91], internal_0n[92]);
  NR2 I105 (internal_0n[100], internal_0n[93], internal_0n[94]);
  NR3 I106 (internal_0n[101], internal_0n[95], internal_0n[96], internal_0n[97]);
  ND4 I107 (out_0d[5], internal_0n[98], internal_0n[99], internal_0n[100], internal_0n[101]);
  ND4 I108 (internal_0n[102], nwayMuxOut_0n[6], nwayMuxOut_1n[6], nwayMuxOut_2n[6], nwayMuxOut_3n[6]);
  ND4 I109 (internal_0n[103], nwayMuxOut_4n[6], nwayMuxOut_5n[6], nwayMuxOut_6n[6], nwayMuxOut_7n[6]);
  ND4 I110 (internal_0n[104], nwayMuxOut_8n[6], nwayMuxOut_9n[6], nwayMuxOut_10n[6], nwayMuxOut_11n[6]);
  ND4 I111 (internal_0n[105], nwayMuxOut_12n[6], nwayMuxOut_13n[6], nwayMuxOut_14n[6], nwayMuxOut_15n[6]);
  ND4 I112 (internal_0n[106], nwayMuxOut_16n[6], nwayMuxOut_17n[6], nwayMuxOut_18n[6], nwayMuxOut_19n[6]);
  ND4 I113 (internal_0n[107], nwayMuxOut_20n[6], nwayMuxOut_21n[6], nwayMuxOut_22n[6], nwayMuxOut_23n[6]);
  ND4 I114 (internal_0n[108], nwayMuxOut_24n[6], nwayMuxOut_25n[6], nwayMuxOut_26n[6], nwayMuxOut_27n[6]);
  ND4 I115 (internal_0n[109], nwayMuxOut_28n[6], nwayMuxOut_29n[6], nwayMuxOut_30n[6], nwayMuxOut_31n[6]);
  ND4 I116 (internal_0n[110], nwayMuxOut_32n[6], nwayMuxOut_33n[6], nwayMuxOut_34n[6], nwayMuxOut_35n[6]);
  ND4 I117 (internal_0n[111], nwayMuxOut_36n[6], nwayMuxOut_37n[6], nwayMuxOut_38n[6], nwayMuxOut_39n[6]);
  ND4 I118 (internal_0n[112], nwayMuxOut_40n[6], nwayMuxOut_41n[6], nwayMuxOut_42n[6], nwayMuxOut_43n[6]);
  ND2 I119 (internal_0n[113], nwayMuxOut_44n[6], nwayMuxOut_45n[6]);
  ND3 I120 (internal_0n[114], nwayMuxOut_46n[6], nwayMuxOut_47n[6], nwayMuxOut_48n[6]);
  NR4 I121 (internal_0n[115], internal_0n[102], internal_0n[103], internal_0n[104], internal_0n[105]);
  NR4 I122 (internal_0n[116], internal_0n[106], internal_0n[107], internal_0n[108], internal_0n[109]);
  NR2 I123 (internal_0n[117], internal_0n[110], internal_0n[111]);
  NR3 I124 (internal_0n[118], internal_0n[112], internal_0n[113], internal_0n[114]);
  ND4 I125 (out_0d[6], internal_0n[115], internal_0n[116], internal_0n[117], internal_0n[118]);
  ND4 I126 (internal_0n[119], nwayMuxOut_0n[7], nwayMuxOut_1n[7], nwayMuxOut_2n[7], nwayMuxOut_3n[7]);
  ND4 I127 (internal_0n[120], nwayMuxOut_4n[7], nwayMuxOut_5n[7], nwayMuxOut_6n[7], nwayMuxOut_7n[7]);
  ND4 I128 (internal_0n[121], nwayMuxOut_8n[7], nwayMuxOut_9n[7], nwayMuxOut_10n[7], nwayMuxOut_11n[7]);
  ND4 I129 (internal_0n[122], nwayMuxOut_12n[7], nwayMuxOut_13n[7], nwayMuxOut_14n[7], nwayMuxOut_15n[7]);
  ND4 I130 (internal_0n[123], nwayMuxOut_16n[7], nwayMuxOut_17n[7], nwayMuxOut_18n[7], nwayMuxOut_19n[7]);
  ND4 I131 (internal_0n[124], nwayMuxOut_20n[7], nwayMuxOut_21n[7], nwayMuxOut_22n[7], nwayMuxOut_23n[7]);
  ND4 I132 (internal_0n[125], nwayMuxOut_24n[7], nwayMuxOut_25n[7], nwayMuxOut_26n[7], nwayMuxOut_27n[7]);
  ND4 I133 (internal_0n[126], nwayMuxOut_28n[7], nwayMuxOut_29n[7], nwayMuxOut_30n[7], nwayMuxOut_31n[7]);
  ND4 I134 (internal_0n[127], nwayMuxOut_32n[7], nwayMuxOut_33n[7], nwayMuxOut_34n[7], nwayMuxOut_35n[7]);
  ND4 I135 (internal_0n[128], nwayMuxOut_36n[7], nwayMuxOut_37n[7], nwayMuxOut_38n[7], nwayMuxOut_39n[7]);
  ND4 I136 (internal_0n[129], nwayMuxOut_40n[7], nwayMuxOut_41n[7], nwayMuxOut_42n[7], nwayMuxOut_43n[7]);
  ND2 I137 (internal_0n[130], nwayMuxOut_44n[7], nwayMuxOut_45n[7]);
  ND3 I138 (internal_0n[131], nwayMuxOut_46n[7], nwayMuxOut_47n[7], nwayMuxOut_48n[7]);
  NR4 I139 (internal_0n[132], internal_0n[119], internal_0n[120], internal_0n[121], internal_0n[122]);
  NR4 I140 (internal_0n[133], internal_0n[123], internal_0n[124], internal_0n[125], internal_0n[126]);
  NR2 I141 (internal_0n[134], internal_0n[127], internal_0n[128]);
  NR3 I142 (internal_0n[135], internal_0n[129], internal_0n[130], internal_0n[131]);
  ND4 I143 (out_0d[7], internal_0n[132], internal_0n[133], internal_0n[134], internal_0n[135]);
  ND4 I144 (internal_0n[136], nwayMuxOut_0n[8], nwayMuxOut_1n[8], nwayMuxOut_2n[8], nwayMuxOut_3n[8]);
  ND4 I145 (internal_0n[137], nwayMuxOut_4n[8], nwayMuxOut_5n[8], nwayMuxOut_6n[8], nwayMuxOut_7n[8]);
  ND4 I146 (internal_0n[138], nwayMuxOut_8n[8], nwayMuxOut_9n[8], nwayMuxOut_10n[8], nwayMuxOut_11n[8]);
  ND4 I147 (internal_0n[139], nwayMuxOut_12n[8], nwayMuxOut_13n[8], nwayMuxOut_14n[8], nwayMuxOut_15n[8]);
  ND4 I148 (internal_0n[140], nwayMuxOut_16n[8], nwayMuxOut_17n[8], nwayMuxOut_18n[8], nwayMuxOut_19n[8]);
  ND4 I149 (internal_0n[141], nwayMuxOut_20n[8], nwayMuxOut_21n[8], nwayMuxOut_22n[8], nwayMuxOut_23n[8]);
  ND4 I150 (internal_0n[142], nwayMuxOut_24n[8], nwayMuxOut_25n[8], nwayMuxOut_26n[8], nwayMuxOut_27n[8]);
  ND4 I151 (internal_0n[143], nwayMuxOut_28n[8], nwayMuxOut_29n[8], nwayMuxOut_30n[8], nwayMuxOut_31n[8]);
  ND4 I152 (internal_0n[144], nwayMuxOut_32n[8], nwayMuxOut_33n[8], nwayMuxOut_34n[8], nwayMuxOut_35n[8]);
  ND4 I153 (internal_0n[145], nwayMuxOut_36n[8], nwayMuxOut_37n[8], nwayMuxOut_38n[8], nwayMuxOut_39n[8]);
  ND4 I154 (internal_0n[146], nwayMuxOut_40n[8], nwayMuxOut_41n[8], nwayMuxOut_42n[8], nwayMuxOut_43n[8]);
  ND2 I155 (internal_0n[147], nwayMuxOut_44n[8], nwayMuxOut_45n[8]);
  ND3 I156 (internal_0n[148], nwayMuxOut_46n[8], nwayMuxOut_47n[8], nwayMuxOut_48n[8]);
  NR4 I157 (internal_0n[149], internal_0n[136], internal_0n[137], internal_0n[138], internal_0n[139]);
  NR4 I158 (internal_0n[150], internal_0n[140], internal_0n[141], internal_0n[142], internal_0n[143]);
  NR2 I159 (internal_0n[151], internal_0n[144], internal_0n[145]);
  NR3 I160 (internal_0n[152], internal_0n[146], internal_0n[147], internal_0n[148]);
  ND4 I161 (out_0d[8], internal_0n[149], internal_0n[150], internal_0n[151], internal_0n[152]);
  ND4 I162 (internal_0n[153], nwayMuxOut_0n[9], nwayMuxOut_1n[9], nwayMuxOut_2n[9], nwayMuxOut_3n[9]);
  ND4 I163 (internal_0n[154], nwayMuxOut_4n[9], nwayMuxOut_5n[9], nwayMuxOut_6n[9], nwayMuxOut_7n[9]);
  ND4 I164 (internal_0n[155], nwayMuxOut_8n[9], nwayMuxOut_9n[9], nwayMuxOut_10n[9], nwayMuxOut_11n[9]);
  ND4 I165 (internal_0n[156], nwayMuxOut_12n[9], nwayMuxOut_13n[9], nwayMuxOut_14n[9], nwayMuxOut_15n[9]);
  ND4 I166 (internal_0n[157], nwayMuxOut_16n[9], nwayMuxOut_17n[9], nwayMuxOut_18n[9], nwayMuxOut_19n[9]);
  ND4 I167 (internal_0n[158], nwayMuxOut_20n[9], nwayMuxOut_21n[9], nwayMuxOut_22n[9], nwayMuxOut_23n[9]);
  ND4 I168 (internal_0n[159], nwayMuxOut_24n[9], nwayMuxOut_25n[9], nwayMuxOut_26n[9], nwayMuxOut_27n[9]);
  ND4 I169 (internal_0n[160], nwayMuxOut_28n[9], nwayMuxOut_29n[9], nwayMuxOut_30n[9], nwayMuxOut_31n[9]);
  ND4 I170 (internal_0n[161], nwayMuxOut_32n[9], nwayMuxOut_33n[9], nwayMuxOut_34n[9], nwayMuxOut_35n[9]);
  ND4 I171 (internal_0n[162], nwayMuxOut_36n[9], nwayMuxOut_37n[9], nwayMuxOut_38n[9], nwayMuxOut_39n[9]);
  ND4 I172 (internal_0n[163], nwayMuxOut_40n[9], nwayMuxOut_41n[9], nwayMuxOut_42n[9], nwayMuxOut_43n[9]);
  ND2 I173 (internal_0n[164], nwayMuxOut_44n[9], nwayMuxOut_45n[9]);
  ND3 I174 (internal_0n[165], nwayMuxOut_46n[9], nwayMuxOut_47n[9], nwayMuxOut_48n[9]);
  NR4 I175 (internal_0n[166], internal_0n[153], internal_0n[154], internal_0n[155], internal_0n[156]);
  NR4 I176 (internal_0n[167], internal_0n[157], internal_0n[158], internal_0n[159], internal_0n[160]);
  NR2 I177 (internal_0n[168], internal_0n[161], internal_0n[162]);
  NR3 I178 (internal_0n[169], internal_0n[163], internal_0n[164], internal_0n[165]);
  ND4 I179 (out_0d[9], internal_0n[166], internal_0n[167], internal_0n[168], internal_0n[169]);
  ND4 I180 (internal_0n[170], nwayMuxOut_0n[10], nwayMuxOut_1n[10], nwayMuxOut_2n[10], nwayMuxOut_3n[10]);
  ND4 I181 (internal_0n[171], nwayMuxOut_4n[10], nwayMuxOut_5n[10], nwayMuxOut_6n[10], nwayMuxOut_7n[10]);
  ND4 I182 (internal_0n[172], nwayMuxOut_8n[10], nwayMuxOut_9n[10], nwayMuxOut_10n[10], nwayMuxOut_11n[10]);
  ND4 I183 (internal_0n[173], nwayMuxOut_12n[10], nwayMuxOut_13n[10], nwayMuxOut_14n[10], nwayMuxOut_15n[10]);
  ND4 I184 (internal_0n[174], nwayMuxOut_16n[10], nwayMuxOut_17n[10], nwayMuxOut_18n[10], nwayMuxOut_19n[10]);
  ND4 I185 (internal_0n[175], nwayMuxOut_20n[10], nwayMuxOut_21n[10], nwayMuxOut_22n[10], nwayMuxOut_23n[10]);
  ND4 I186 (internal_0n[176], nwayMuxOut_24n[10], nwayMuxOut_25n[10], nwayMuxOut_26n[10], nwayMuxOut_27n[10]);
  ND4 I187 (internal_0n[177], nwayMuxOut_28n[10], nwayMuxOut_29n[10], nwayMuxOut_30n[10], nwayMuxOut_31n[10]);
  ND4 I188 (internal_0n[178], nwayMuxOut_32n[10], nwayMuxOut_33n[10], nwayMuxOut_34n[10], nwayMuxOut_35n[10]);
  ND4 I189 (internal_0n[179], nwayMuxOut_36n[10], nwayMuxOut_37n[10], nwayMuxOut_38n[10], nwayMuxOut_39n[10]);
  ND4 I190 (internal_0n[180], nwayMuxOut_40n[10], nwayMuxOut_41n[10], nwayMuxOut_42n[10], nwayMuxOut_43n[10]);
  ND2 I191 (internal_0n[181], nwayMuxOut_44n[10], nwayMuxOut_45n[10]);
  ND3 I192 (internal_0n[182], nwayMuxOut_46n[10], nwayMuxOut_47n[10], nwayMuxOut_48n[10]);
  NR4 I193 (internal_0n[183], internal_0n[170], internal_0n[171], internal_0n[172], internal_0n[173]);
  NR4 I194 (internal_0n[184], internal_0n[174], internal_0n[175], internal_0n[176], internal_0n[177]);
  NR2 I195 (internal_0n[185], internal_0n[178], internal_0n[179]);
  NR3 I196 (internal_0n[186], internal_0n[180], internal_0n[181], internal_0n[182]);
  ND4 I197 (out_0d[10], internal_0n[183], internal_0n[184], internal_0n[185], internal_0n[186]);
  ND4 I198 (internal_0n[187], nwayMuxOut_0n[11], nwayMuxOut_1n[11], nwayMuxOut_2n[11], nwayMuxOut_3n[11]);
  ND4 I199 (internal_0n[188], nwayMuxOut_4n[11], nwayMuxOut_5n[11], nwayMuxOut_6n[11], nwayMuxOut_7n[11]);
  ND4 I200 (internal_0n[189], nwayMuxOut_8n[11], nwayMuxOut_9n[11], nwayMuxOut_10n[11], nwayMuxOut_11n[11]);
  ND4 I201 (internal_0n[190], nwayMuxOut_12n[11], nwayMuxOut_13n[11], nwayMuxOut_14n[11], nwayMuxOut_15n[11]);
  ND4 I202 (internal_0n[191], nwayMuxOut_16n[11], nwayMuxOut_17n[11], nwayMuxOut_18n[11], nwayMuxOut_19n[11]);
  ND4 I203 (internal_0n[192], nwayMuxOut_20n[11], nwayMuxOut_21n[11], nwayMuxOut_22n[11], nwayMuxOut_23n[11]);
  ND4 I204 (internal_0n[193], nwayMuxOut_24n[11], nwayMuxOut_25n[11], nwayMuxOut_26n[11], nwayMuxOut_27n[11]);
  ND4 I205 (internal_0n[194], nwayMuxOut_28n[11], nwayMuxOut_29n[11], nwayMuxOut_30n[11], nwayMuxOut_31n[11]);
  ND4 I206 (internal_0n[195], nwayMuxOut_32n[11], nwayMuxOut_33n[11], nwayMuxOut_34n[11], nwayMuxOut_35n[11]);
  ND4 I207 (internal_0n[196], nwayMuxOut_36n[11], nwayMuxOut_37n[11], nwayMuxOut_38n[11], nwayMuxOut_39n[11]);
  ND4 I208 (internal_0n[197], nwayMuxOut_40n[11], nwayMuxOut_41n[11], nwayMuxOut_42n[11], nwayMuxOut_43n[11]);
  ND2 I209 (internal_0n[198], nwayMuxOut_44n[11], nwayMuxOut_45n[11]);
  ND3 I210 (internal_0n[199], nwayMuxOut_46n[11], nwayMuxOut_47n[11], nwayMuxOut_48n[11]);
  NR4 I211 (internal_0n[200], internal_0n[187], internal_0n[188], internal_0n[189], internal_0n[190]);
  NR4 I212 (internal_0n[201], internal_0n[191], internal_0n[192], internal_0n[193], internal_0n[194]);
  NR2 I213 (internal_0n[202], internal_0n[195], internal_0n[196]);
  NR3 I214 (internal_0n[203], internal_0n[197], internal_0n[198], internal_0n[199]);
  ND4 I215 (out_0d[11], internal_0n[200], internal_0n[201], internal_0n[202], internal_0n[203]);
  ND4 I216 (internal_0n[204], nwayMuxOut_0n[12], nwayMuxOut_1n[12], nwayMuxOut_2n[12], nwayMuxOut_3n[12]);
  ND4 I217 (internal_0n[205], nwayMuxOut_4n[12], nwayMuxOut_5n[12], nwayMuxOut_6n[12], nwayMuxOut_7n[12]);
  ND4 I218 (internal_0n[206], nwayMuxOut_8n[12], nwayMuxOut_9n[12], nwayMuxOut_10n[12], nwayMuxOut_11n[12]);
  ND4 I219 (internal_0n[207], nwayMuxOut_12n[12], nwayMuxOut_13n[12], nwayMuxOut_14n[12], nwayMuxOut_15n[12]);
  ND4 I220 (internal_0n[208], nwayMuxOut_16n[12], nwayMuxOut_17n[12], nwayMuxOut_18n[12], nwayMuxOut_19n[12]);
  ND4 I221 (internal_0n[209], nwayMuxOut_20n[12], nwayMuxOut_21n[12], nwayMuxOut_22n[12], nwayMuxOut_23n[12]);
  ND4 I222 (internal_0n[210], nwayMuxOut_24n[12], nwayMuxOut_25n[12], nwayMuxOut_26n[12], nwayMuxOut_27n[12]);
  ND4 I223 (internal_0n[211], nwayMuxOut_28n[12], nwayMuxOut_29n[12], nwayMuxOut_30n[12], nwayMuxOut_31n[12]);
  ND4 I224 (internal_0n[212], nwayMuxOut_32n[12], nwayMuxOut_33n[12], nwayMuxOut_34n[12], nwayMuxOut_35n[12]);
  ND4 I225 (internal_0n[213], nwayMuxOut_36n[12], nwayMuxOut_37n[12], nwayMuxOut_38n[12], nwayMuxOut_39n[12]);
  ND4 I226 (internal_0n[214], nwayMuxOut_40n[12], nwayMuxOut_41n[12], nwayMuxOut_42n[12], nwayMuxOut_43n[12]);
  ND2 I227 (internal_0n[215], nwayMuxOut_44n[12], nwayMuxOut_45n[12]);
  ND3 I228 (internal_0n[216], nwayMuxOut_46n[12], nwayMuxOut_47n[12], nwayMuxOut_48n[12]);
  NR4 I229 (internal_0n[217], internal_0n[204], internal_0n[205], internal_0n[206], internal_0n[207]);
  NR4 I230 (internal_0n[218], internal_0n[208], internal_0n[209], internal_0n[210], internal_0n[211]);
  NR2 I231 (internal_0n[219], internal_0n[212], internal_0n[213]);
  NR3 I232 (internal_0n[220], internal_0n[214], internal_0n[215], internal_0n[216]);
  ND4 I233 (out_0d[12], internal_0n[217], internal_0n[218], internal_0n[219], internal_0n[220]);
  ND4 I234 (internal_0n[221], nwayMuxOut_0n[13], nwayMuxOut_1n[13], nwayMuxOut_2n[13], nwayMuxOut_3n[13]);
  ND4 I235 (internal_0n[222], nwayMuxOut_4n[13], nwayMuxOut_5n[13], nwayMuxOut_6n[13], nwayMuxOut_7n[13]);
  ND4 I236 (internal_0n[223], nwayMuxOut_8n[13], nwayMuxOut_9n[13], nwayMuxOut_10n[13], nwayMuxOut_11n[13]);
  ND4 I237 (internal_0n[224], nwayMuxOut_12n[13], nwayMuxOut_13n[13], nwayMuxOut_14n[13], nwayMuxOut_15n[13]);
  ND4 I238 (internal_0n[225], nwayMuxOut_16n[13], nwayMuxOut_17n[13], nwayMuxOut_18n[13], nwayMuxOut_19n[13]);
  ND4 I239 (internal_0n[226], nwayMuxOut_20n[13], nwayMuxOut_21n[13], nwayMuxOut_22n[13], nwayMuxOut_23n[13]);
  ND4 I240 (internal_0n[227], nwayMuxOut_24n[13], nwayMuxOut_25n[13], nwayMuxOut_26n[13], nwayMuxOut_27n[13]);
  ND4 I241 (internal_0n[228], nwayMuxOut_28n[13], nwayMuxOut_29n[13], nwayMuxOut_30n[13], nwayMuxOut_31n[13]);
  ND4 I242 (internal_0n[229], nwayMuxOut_32n[13], nwayMuxOut_33n[13], nwayMuxOut_34n[13], nwayMuxOut_35n[13]);
  ND4 I243 (internal_0n[230], nwayMuxOut_36n[13], nwayMuxOut_37n[13], nwayMuxOut_38n[13], nwayMuxOut_39n[13]);
  ND4 I244 (internal_0n[231], nwayMuxOut_40n[13], nwayMuxOut_41n[13], nwayMuxOut_42n[13], nwayMuxOut_43n[13]);
  ND2 I245 (internal_0n[232], nwayMuxOut_44n[13], nwayMuxOut_45n[13]);
  ND3 I246 (internal_0n[233], nwayMuxOut_46n[13], nwayMuxOut_47n[13], nwayMuxOut_48n[13]);
  NR4 I247 (internal_0n[234], internal_0n[221], internal_0n[222], internal_0n[223], internal_0n[224]);
  NR4 I248 (internal_0n[235], internal_0n[225], internal_0n[226], internal_0n[227], internal_0n[228]);
  NR2 I249 (internal_0n[236], internal_0n[229], internal_0n[230]);
  NR3 I250 (internal_0n[237], internal_0n[231], internal_0n[232], internal_0n[233]);
  ND4 I251 (out_0d[13], internal_0n[234], internal_0n[235], internal_0n[236], internal_0n[237]);
  ND4 I252 (internal_0n[238], nwayMuxOut_0n[14], nwayMuxOut_1n[14], nwayMuxOut_2n[14], nwayMuxOut_3n[14]);
  ND4 I253 (internal_0n[239], nwayMuxOut_4n[14], nwayMuxOut_5n[14], nwayMuxOut_6n[14], nwayMuxOut_7n[14]);
  ND4 I254 (internal_0n[240], nwayMuxOut_8n[14], nwayMuxOut_9n[14], nwayMuxOut_10n[14], nwayMuxOut_11n[14]);
  ND4 I255 (internal_0n[241], nwayMuxOut_12n[14], nwayMuxOut_13n[14], nwayMuxOut_14n[14], nwayMuxOut_15n[14]);
  ND4 I256 (internal_0n[242], nwayMuxOut_16n[14], nwayMuxOut_17n[14], nwayMuxOut_18n[14], nwayMuxOut_19n[14]);
  ND4 I257 (internal_0n[243], nwayMuxOut_20n[14], nwayMuxOut_21n[14], nwayMuxOut_22n[14], nwayMuxOut_23n[14]);
  ND4 I258 (internal_0n[244], nwayMuxOut_24n[14], nwayMuxOut_25n[14], nwayMuxOut_26n[14], nwayMuxOut_27n[14]);
  ND4 I259 (internal_0n[245], nwayMuxOut_28n[14], nwayMuxOut_29n[14], nwayMuxOut_30n[14], nwayMuxOut_31n[14]);
  ND4 I260 (internal_0n[246], nwayMuxOut_32n[14], nwayMuxOut_33n[14], nwayMuxOut_34n[14], nwayMuxOut_35n[14]);
  ND4 I261 (internal_0n[247], nwayMuxOut_36n[14], nwayMuxOut_37n[14], nwayMuxOut_38n[14], nwayMuxOut_39n[14]);
  ND4 I262 (internal_0n[248], nwayMuxOut_40n[14], nwayMuxOut_41n[14], nwayMuxOut_42n[14], nwayMuxOut_43n[14]);
  ND2 I263 (internal_0n[249], nwayMuxOut_44n[14], nwayMuxOut_45n[14]);
  ND3 I264 (internal_0n[250], nwayMuxOut_46n[14], nwayMuxOut_47n[14], nwayMuxOut_48n[14]);
  NR4 I265 (internal_0n[251], internal_0n[238], internal_0n[239], internal_0n[240], internal_0n[241]);
  NR4 I266 (internal_0n[252], internal_0n[242], internal_0n[243], internal_0n[244], internal_0n[245]);
  NR2 I267 (internal_0n[253], internal_0n[246], internal_0n[247]);
  NR3 I268 (internal_0n[254], internal_0n[248], internal_0n[249], internal_0n[250]);
  ND4 I269 (out_0d[14], internal_0n[251], internal_0n[252], internal_0n[253], internal_0n[254]);
  ND4 I270 (internal_0n[255], nwayMuxOut_0n[15], nwayMuxOut_1n[15], nwayMuxOut_2n[15], nwayMuxOut_3n[15]);
  ND4 I271 (internal_0n[256], nwayMuxOut_4n[15], nwayMuxOut_5n[15], nwayMuxOut_6n[15], nwayMuxOut_7n[15]);
  ND4 I272 (internal_0n[257], nwayMuxOut_8n[15], nwayMuxOut_9n[15], nwayMuxOut_10n[15], nwayMuxOut_11n[15]);
  ND4 I273 (internal_0n[258], nwayMuxOut_12n[15], nwayMuxOut_13n[15], nwayMuxOut_14n[15], nwayMuxOut_15n[15]);
  ND4 I274 (internal_0n[259], nwayMuxOut_16n[15], nwayMuxOut_17n[15], nwayMuxOut_18n[15], nwayMuxOut_19n[15]);
  ND4 I275 (internal_0n[260], nwayMuxOut_20n[15], nwayMuxOut_21n[15], nwayMuxOut_22n[15], nwayMuxOut_23n[15]);
  ND4 I276 (internal_0n[261], nwayMuxOut_24n[15], nwayMuxOut_25n[15], nwayMuxOut_26n[15], nwayMuxOut_27n[15]);
  ND4 I277 (internal_0n[262], nwayMuxOut_28n[15], nwayMuxOut_29n[15], nwayMuxOut_30n[15], nwayMuxOut_31n[15]);
  ND4 I278 (internal_0n[263], nwayMuxOut_32n[15], nwayMuxOut_33n[15], nwayMuxOut_34n[15], nwayMuxOut_35n[15]);
  ND4 I279 (internal_0n[264], nwayMuxOut_36n[15], nwayMuxOut_37n[15], nwayMuxOut_38n[15], nwayMuxOut_39n[15]);
  ND4 I280 (internal_0n[265], nwayMuxOut_40n[15], nwayMuxOut_41n[15], nwayMuxOut_42n[15], nwayMuxOut_43n[15]);
  ND2 I281 (internal_0n[266], nwayMuxOut_44n[15], nwayMuxOut_45n[15]);
  ND3 I282 (internal_0n[267], nwayMuxOut_46n[15], nwayMuxOut_47n[15], nwayMuxOut_48n[15]);
  NR4 I283 (internal_0n[268], internal_0n[255], internal_0n[256], internal_0n[257], internal_0n[258]);
  NR4 I284 (internal_0n[269], internal_0n[259], internal_0n[260], internal_0n[261], internal_0n[262]);
  NR2 I285 (internal_0n[270], internal_0n[263], internal_0n[264]);
  NR3 I286 (internal_0n[271], internal_0n[265], internal_0n[266], internal_0n[267]);
  ND4 I287 (out_0d[15], internal_0n[268], internal_0n[269], internal_0n[270], internal_0n[271]);
  ND4 I288 (internal_0n[272], nwayMuxOut_0n[16], nwayMuxOut_1n[16], nwayMuxOut_2n[16], nwayMuxOut_3n[16]);
  ND4 I289 (internal_0n[273], nwayMuxOut_4n[16], nwayMuxOut_5n[16], nwayMuxOut_6n[16], nwayMuxOut_7n[16]);
  ND4 I290 (internal_0n[274], nwayMuxOut_8n[16], nwayMuxOut_9n[16], nwayMuxOut_10n[16], nwayMuxOut_11n[16]);
  ND4 I291 (internal_0n[275], nwayMuxOut_12n[16], nwayMuxOut_13n[16], nwayMuxOut_14n[16], nwayMuxOut_15n[16]);
  ND4 I292 (internal_0n[276], nwayMuxOut_16n[16], nwayMuxOut_17n[16], nwayMuxOut_18n[16], nwayMuxOut_19n[16]);
  ND4 I293 (internal_0n[277], nwayMuxOut_20n[16], nwayMuxOut_21n[16], nwayMuxOut_22n[16], nwayMuxOut_23n[16]);
  ND4 I294 (internal_0n[278], nwayMuxOut_24n[16], nwayMuxOut_25n[16], nwayMuxOut_26n[16], nwayMuxOut_27n[16]);
  ND4 I295 (internal_0n[279], nwayMuxOut_28n[16], nwayMuxOut_29n[16], nwayMuxOut_30n[16], nwayMuxOut_31n[16]);
  ND4 I296 (internal_0n[280], nwayMuxOut_32n[16], nwayMuxOut_33n[16], nwayMuxOut_34n[16], nwayMuxOut_35n[16]);
  ND4 I297 (internal_0n[281], nwayMuxOut_36n[16], nwayMuxOut_37n[16], nwayMuxOut_38n[16], nwayMuxOut_39n[16]);
  ND4 I298 (internal_0n[282], nwayMuxOut_40n[16], nwayMuxOut_41n[16], nwayMuxOut_42n[16], nwayMuxOut_43n[16]);
  ND2 I299 (internal_0n[283], nwayMuxOut_44n[16], nwayMuxOut_45n[16]);
  ND3 I300 (internal_0n[284], nwayMuxOut_46n[16], nwayMuxOut_47n[16], nwayMuxOut_48n[16]);
  NR4 I301 (internal_0n[285], internal_0n[272], internal_0n[273], internal_0n[274], internal_0n[275]);
  NR4 I302 (internal_0n[286], internal_0n[276], internal_0n[277], internal_0n[278], internal_0n[279]);
  NR2 I303 (internal_0n[287], internal_0n[280], internal_0n[281]);
  NR3 I304 (internal_0n[288], internal_0n[282], internal_0n[283], internal_0n[284]);
  ND4 I305 (out_0d[16], internal_0n[285], internal_0n[286], internal_0n[287], internal_0n[288]);
  ND4 I306 (internal_0n[289], nwayMuxOut_0n[17], nwayMuxOut_1n[17], nwayMuxOut_2n[17], nwayMuxOut_3n[17]);
  ND4 I307 (internal_0n[290], nwayMuxOut_4n[17], nwayMuxOut_5n[17], nwayMuxOut_6n[17], nwayMuxOut_7n[17]);
  ND4 I308 (internal_0n[291], nwayMuxOut_8n[17], nwayMuxOut_9n[17], nwayMuxOut_10n[17], nwayMuxOut_11n[17]);
  ND4 I309 (internal_0n[292], nwayMuxOut_12n[17], nwayMuxOut_13n[17], nwayMuxOut_14n[17], nwayMuxOut_15n[17]);
  ND4 I310 (internal_0n[293], nwayMuxOut_16n[17], nwayMuxOut_17n[17], nwayMuxOut_18n[17], nwayMuxOut_19n[17]);
  ND4 I311 (internal_0n[294], nwayMuxOut_20n[17], nwayMuxOut_21n[17], nwayMuxOut_22n[17], nwayMuxOut_23n[17]);
  ND4 I312 (internal_0n[295], nwayMuxOut_24n[17], nwayMuxOut_25n[17], nwayMuxOut_26n[17], nwayMuxOut_27n[17]);
  ND4 I313 (internal_0n[296], nwayMuxOut_28n[17], nwayMuxOut_29n[17], nwayMuxOut_30n[17], nwayMuxOut_31n[17]);
  ND4 I314 (internal_0n[297], nwayMuxOut_32n[17], nwayMuxOut_33n[17], nwayMuxOut_34n[17], nwayMuxOut_35n[17]);
  ND4 I315 (internal_0n[298], nwayMuxOut_36n[17], nwayMuxOut_37n[17], nwayMuxOut_38n[17], nwayMuxOut_39n[17]);
  ND4 I316 (internal_0n[299], nwayMuxOut_40n[17], nwayMuxOut_41n[17], nwayMuxOut_42n[17], nwayMuxOut_43n[17]);
  ND2 I317 (internal_0n[300], nwayMuxOut_44n[17], nwayMuxOut_45n[17]);
  ND3 I318 (internal_0n[301], nwayMuxOut_46n[17], nwayMuxOut_47n[17], nwayMuxOut_48n[17]);
  NR4 I319 (internal_0n[302], internal_0n[289], internal_0n[290], internal_0n[291], internal_0n[292]);
  NR4 I320 (internal_0n[303], internal_0n[293], internal_0n[294], internal_0n[295], internal_0n[296]);
  NR2 I321 (internal_0n[304], internal_0n[297], internal_0n[298]);
  NR3 I322 (internal_0n[305], internal_0n[299], internal_0n[300], internal_0n[301]);
  ND4 I323 (out_0d[17], internal_0n[302], internal_0n[303], internal_0n[304], internal_0n[305]);
  ND4 I324 (internal_0n[306], nwayMuxOut_0n[18], nwayMuxOut_1n[18], nwayMuxOut_2n[18], nwayMuxOut_3n[18]);
  ND4 I325 (internal_0n[307], nwayMuxOut_4n[18], nwayMuxOut_5n[18], nwayMuxOut_6n[18], nwayMuxOut_7n[18]);
  ND4 I326 (internal_0n[308], nwayMuxOut_8n[18], nwayMuxOut_9n[18], nwayMuxOut_10n[18], nwayMuxOut_11n[18]);
  ND4 I327 (internal_0n[309], nwayMuxOut_12n[18], nwayMuxOut_13n[18], nwayMuxOut_14n[18], nwayMuxOut_15n[18]);
  ND4 I328 (internal_0n[310], nwayMuxOut_16n[18], nwayMuxOut_17n[18], nwayMuxOut_18n[18], nwayMuxOut_19n[18]);
  ND4 I329 (internal_0n[311], nwayMuxOut_20n[18], nwayMuxOut_21n[18], nwayMuxOut_22n[18], nwayMuxOut_23n[18]);
  ND4 I330 (internal_0n[312], nwayMuxOut_24n[18], nwayMuxOut_25n[18], nwayMuxOut_26n[18], nwayMuxOut_27n[18]);
  ND4 I331 (internal_0n[313], nwayMuxOut_28n[18], nwayMuxOut_29n[18], nwayMuxOut_30n[18], nwayMuxOut_31n[18]);
  ND4 I332 (internal_0n[314], nwayMuxOut_32n[18], nwayMuxOut_33n[18], nwayMuxOut_34n[18], nwayMuxOut_35n[18]);
  ND4 I333 (internal_0n[315], nwayMuxOut_36n[18], nwayMuxOut_37n[18], nwayMuxOut_38n[18], nwayMuxOut_39n[18]);
  ND4 I334 (internal_0n[316], nwayMuxOut_40n[18], nwayMuxOut_41n[18], nwayMuxOut_42n[18], nwayMuxOut_43n[18]);
  ND2 I335 (internal_0n[317], nwayMuxOut_44n[18], nwayMuxOut_45n[18]);
  ND3 I336 (internal_0n[318], nwayMuxOut_46n[18], nwayMuxOut_47n[18], nwayMuxOut_48n[18]);
  NR4 I337 (internal_0n[319], internal_0n[306], internal_0n[307], internal_0n[308], internal_0n[309]);
  NR4 I338 (internal_0n[320], internal_0n[310], internal_0n[311], internal_0n[312], internal_0n[313]);
  NR2 I339 (internal_0n[321], internal_0n[314], internal_0n[315]);
  NR3 I340 (internal_0n[322], internal_0n[316], internal_0n[317], internal_0n[318]);
  ND4 I341 (out_0d[18], internal_0n[319], internal_0n[320], internal_0n[321], internal_0n[322]);
  ND4 I342 (internal_0n[323], nwayMuxOut_0n[19], nwayMuxOut_1n[19], nwayMuxOut_2n[19], nwayMuxOut_3n[19]);
  ND4 I343 (internal_0n[324], nwayMuxOut_4n[19], nwayMuxOut_5n[19], nwayMuxOut_6n[19], nwayMuxOut_7n[19]);
  ND4 I344 (internal_0n[325], nwayMuxOut_8n[19], nwayMuxOut_9n[19], nwayMuxOut_10n[19], nwayMuxOut_11n[19]);
  ND4 I345 (internal_0n[326], nwayMuxOut_12n[19], nwayMuxOut_13n[19], nwayMuxOut_14n[19], nwayMuxOut_15n[19]);
  ND4 I346 (internal_0n[327], nwayMuxOut_16n[19], nwayMuxOut_17n[19], nwayMuxOut_18n[19], nwayMuxOut_19n[19]);
  ND4 I347 (internal_0n[328], nwayMuxOut_20n[19], nwayMuxOut_21n[19], nwayMuxOut_22n[19], nwayMuxOut_23n[19]);
  ND4 I348 (internal_0n[329], nwayMuxOut_24n[19], nwayMuxOut_25n[19], nwayMuxOut_26n[19], nwayMuxOut_27n[19]);
  ND4 I349 (internal_0n[330], nwayMuxOut_28n[19], nwayMuxOut_29n[19], nwayMuxOut_30n[19], nwayMuxOut_31n[19]);
  ND4 I350 (internal_0n[331], nwayMuxOut_32n[19], nwayMuxOut_33n[19], nwayMuxOut_34n[19], nwayMuxOut_35n[19]);
  ND4 I351 (internal_0n[332], nwayMuxOut_36n[19], nwayMuxOut_37n[19], nwayMuxOut_38n[19], nwayMuxOut_39n[19]);
  ND4 I352 (internal_0n[333], nwayMuxOut_40n[19], nwayMuxOut_41n[19], nwayMuxOut_42n[19], nwayMuxOut_43n[19]);
  ND2 I353 (internal_0n[334], nwayMuxOut_44n[19], nwayMuxOut_45n[19]);
  ND3 I354 (internal_0n[335], nwayMuxOut_46n[19], nwayMuxOut_47n[19], nwayMuxOut_48n[19]);
  NR4 I355 (internal_0n[336], internal_0n[323], internal_0n[324], internal_0n[325], internal_0n[326]);
  NR4 I356 (internal_0n[337], internal_0n[327], internal_0n[328], internal_0n[329], internal_0n[330]);
  NR2 I357 (internal_0n[338], internal_0n[331], internal_0n[332]);
  NR3 I358 (internal_0n[339], internal_0n[333], internal_0n[334], internal_0n[335]);
  ND4 I359 (out_0d[19], internal_0n[336], internal_0n[337], internal_0n[338], internal_0n[339]);
  ND4 I360 (internal_0n[340], nwayMuxOut_0n[20], nwayMuxOut_1n[20], nwayMuxOut_2n[20], nwayMuxOut_3n[20]);
  ND4 I361 (internal_0n[341], nwayMuxOut_4n[20], nwayMuxOut_5n[20], nwayMuxOut_6n[20], nwayMuxOut_7n[20]);
  ND4 I362 (internal_0n[342], nwayMuxOut_8n[20], nwayMuxOut_9n[20], nwayMuxOut_10n[20], nwayMuxOut_11n[20]);
  ND4 I363 (internal_0n[343], nwayMuxOut_12n[20], nwayMuxOut_13n[20], nwayMuxOut_14n[20], nwayMuxOut_15n[20]);
  ND4 I364 (internal_0n[344], nwayMuxOut_16n[20], nwayMuxOut_17n[20], nwayMuxOut_18n[20], nwayMuxOut_19n[20]);
  ND4 I365 (internal_0n[345], nwayMuxOut_20n[20], nwayMuxOut_21n[20], nwayMuxOut_22n[20], nwayMuxOut_23n[20]);
  ND4 I366 (internal_0n[346], nwayMuxOut_24n[20], nwayMuxOut_25n[20], nwayMuxOut_26n[20], nwayMuxOut_27n[20]);
  ND4 I367 (internal_0n[347], nwayMuxOut_28n[20], nwayMuxOut_29n[20], nwayMuxOut_30n[20], nwayMuxOut_31n[20]);
  ND4 I368 (internal_0n[348], nwayMuxOut_32n[20], nwayMuxOut_33n[20], nwayMuxOut_34n[20], nwayMuxOut_35n[20]);
  ND4 I369 (internal_0n[349], nwayMuxOut_36n[20], nwayMuxOut_37n[20], nwayMuxOut_38n[20], nwayMuxOut_39n[20]);
  ND4 I370 (internal_0n[350], nwayMuxOut_40n[20], nwayMuxOut_41n[20], nwayMuxOut_42n[20], nwayMuxOut_43n[20]);
  ND2 I371 (internal_0n[351], nwayMuxOut_44n[20], nwayMuxOut_45n[20]);
  ND3 I372 (internal_0n[352], nwayMuxOut_46n[20], nwayMuxOut_47n[20], nwayMuxOut_48n[20]);
  NR4 I373 (internal_0n[353], internal_0n[340], internal_0n[341], internal_0n[342], internal_0n[343]);
  NR4 I374 (internal_0n[354], internal_0n[344], internal_0n[345], internal_0n[346], internal_0n[347]);
  NR2 I375 (internal_0n[355], internal_0n[348], internal_0n[349]);
  NR3 I376 (internal_0n[356], internal_0n[350], internal_0n[351], internal_0n[352]);
  ND4 I377 (out_0d[20], internal_0n[353], internal_0n[354], internal_0n[355], internal_0n[356]);
  ND4 I378 (internal_0n[357], nwayMuxOut_0n[21], nwayMuxOut_1n[21], nwayMuxOut_2n[21], nwayMuxOut_3n[21]);
  ND4 I379 (internal_0n[358], nwayMuxOut_4n[21], nwayMuxOut_5n[21], nwayMuxOut_6n[21], nwayMuxOut_7n[21]);
  ND4 I380 (internal_0n[359], nwayMuxOut_8n[21], nwayMuxOut_9n[21], nwayMuxOut_10n[21], nwayMuxOut_11n[21]);
  ND4 I381 (internal_0n[360], nwayMuxOut_12n[21], nwayMuxOut_13n[21], nwayMuxOut_14n[21], nwayMuxOut_15n[21]);
  ND4 I382 (internal_0n[361], nwayMuxOut_16n[21], nwayMuxOut_17n[21], nwayMuxOut_18n[21], nwayMuxOut_19n[21]);
  ND4 I383 (internal_0n[362], nwayMuxOut_20n[21], nwayMuxOut_21n[21], nwayMuxOut_22n[21], nwayMuxOut_23n[21]);
  ND4 I384 (internal_0n[363], nwayMuxOut_24n[21], nwayMuxOut_25n[21], nwayMuxOut_26n[21], nwayMuxOut_27n[21]);
  ND4 I385 (internal_0n[364], nwayMuxOut_28n[21], nwayMuxOut_29n[21], nwayMuxOut_30n[21], nwayMuxOut_31n[21]);
  ND4 I386 (internal_0n[365], nwayMuxOut_32n[21], nwayMuxOut_33n[21], nwayMuxOut_34n[21], nwayMuxOut_35n[21]);
  ND4 I387 (internal_0n[366], nwayMuxOut_36n[21], nwayMuxOut_37n[21], nwayMuxOut_38n[21], nwayMuxOut_39n[21]);
  ND4 I388 (internal_0n[367], nwayMuxOut_40n[21], nwayMuxOut_41n[21], nwayMuxOut_42n[21], nwayMuxOut_43n[21]);
  ND2 I389 (internal_0n[368], nwayMuxOut_44n[21], nwayMuxOut_45n[21]);
  ND3 I390 (internal_0n[369], nwayMuxOut_46n[21], nwayMuxOut_47n[21], nwayMuxOut_48n[21]);
  NR4 I391 (internal_0n[370], internal_0n[357], internal_0n[358], internal_0n[359], internal_0n[360]);
  NR4 I392 (internal_0n[371], internal_0n[361], internal_0n[362], internal_0n[363], internal_0n[364]);
  NR2 I393 (internal_0n[372], internal_0n[365], internal_0n[366]);
  NR3 I394 (internal_0n[373], internal_0n[367], internal_0n[368], internal_0n[369]);
  ND4 I395 (out_0d[21], internal_0n[370], internal_0n[371], internal_0n[372], internal_0n[373]);
  ND4 I396 (internal_0n[374], nwayMuxOut_0n[22], nwayMuxOut_1n[22], nwayMuxOut_2n[22], nwayMuxOut_3n[22]);
  ND4 I397 (internal_0n[375], nwayMuxOut_4n[22], nwayMuxOut_5n[22], nwayMuxOut_6n[22], nwayMuxOut_7n[22]);
  ND4 I398 (internal_0n[376], nwayMuxOut_8n[22], nwayMuxOut_9n[22], nwayMuxOut_10n[22], nwayMuxOut_11n[22]);
  ND4 I399 (internal_0n[377], nwayMuxOut_12n[22], nwayMuxOut_13n[22], nwayMuxOut_14n[22], nwayMuxOut_15n[22]);
  ND4 I400 (internal_0n[378], nwayMuxOut_16n[22], nwayMuxOut_17n[22], nwayMuxOut_18n[22], nwayMuxOut_19n[22]);
  ND4 I401 (internal_0n[379], nwayMuxOut_20n[22], nwayMuxOut_21n[22], nwayMuxOut_22n[22], nwayMuxOut_23n[22]);
  ND4 I402 (internal_0n[380], nwayMuxOut_24n[22], nwayMuxOut_25n[22], nwayMuxOut_26n[22], nwayMuxOut_27n[22]);
  ND4 I403 (internal_0n[381], nwayMuxOut_28n[22], nwayMuxOut_29n[22], nwayMuxOut_30n[22], nwayMuxOut_31n[22]);
  ND4 I404 (internal_0n[382], nwayMuxOut_32n[22], nwayMuxOut_33n[22], nwayMuxOut_34n[22], nwayMuxOut_35n[22]);
  ND4 I405 (internal_0n[383], nwayMuxOut_36n[22], nwayMuxOut_37n[22], nwayMuxOut_38n[22], nwayMuxOut_39n[22]);
  ND4 I406 (internal_0n[384], nwayMuxOut_40n[22], nwayMuxOut_41n[22], nwayMuxOut_42n[22], nwayMuxOut_43n[22]);
  ND2 I407 (internal_0n[385], nwayMuxOut_44n[22], nwayMuxOut_45n[22]);
  ND3 I408 (internal_0n[386], nwayMuxOut_46n[22], nwayMuxOut_47n[22], nwayMuxOut_48n[22]);
  NR4 I409 (internal_0n[387], internal_0n[374], internal_0n[375], internal_0n[376], internal_0n[377]);
  NR4 I410 (internal_0n[388], internal_0n[378], internal_0n[379], internal_0n[380], internal_0n[381]);
  NR2 I411 (internal_0n[389], internal_0n[382], internal_0n[383]);
  NR3 I412 (internal_0n[390], internal_0n[384], internal_0n[385], internal_0n[386]);
  ND4 I413 (out_0d[22], internal_0n[387], internal_0n[388], internal_0n[389], internal_0n[390]);
  ND4 I414 (internal_0n[391], nwayMuxOut_0n[23], nwayMuxOut_1n[23], nwayMuxOut_2n[23], nwayMuxOut_3n[23]);
  ND4 I415 (internal_0n[392], nwayMuxOut_4n[23], nwayMuxOut_5n[23], nwayMuxOut_6n[23], nwayMuxOut_7n[23]);
  ND4 I416 (internal_0n[393], nwayMuxOut_8n[23], nwayMuxOut_9n[23], nwayMuxOut_10n[23], nwayMuxOut_11n[23]);
  ND4 I417 (internal_0n[394], nwayMuxOut_12n[23], nwayMuxOut_13n[23], nwayMuxOut_14n[23], nwayMuxOut_15n[23]);
  ND4 I418 (internal_0n[395], nwayMuxOut_16n[23], nwayMuxOut_17n[23], nwayMuxOut_18n[23], nwayMuxOut_19n[23]);
  ND4 I419 (internal_0n[396], nwayMuxOut_20n[23], nwayMuxOut_21n[23], nwayMuxOut_22n[23], nwayMuxOut_23n[23]);
  ND4 I420 (internal_0n[397], nwayMuxOut_24n[23], nwayMuxOut_25n[23], nwayMuxOut_26n[23], nwayMuxOut_27n[23]);
  ND4 I421 (internal_0n[398], nwayMuxOut_28n[23], nwayMuxOut_29n[23], nwayMuxOut_30n[23], nwayMuxOut_31n[23]);
  ND4 I422 (internal_0n[399], nwayMuxOut_32n[23], nwayMuxOut_33n[23], nwayMuxOut_34n[23], nwayMuxOut_35n[23]);
  ND4 I423 (internal_0n[400], nwayMuxOut_36n[23], nwayMuxOut_37n[23], nwayMuxOut_38n[23], nwayMuxOut_39n[23]);
  ND4 I424 (internal_0n[401], nwayMuxOut_40n[23], nwayMuxOut_41n[23], nwayMuxOut_42n[23], nwayMuxOut_43n[23]);
  ND2 I425 (internal_0n[402], nwayMuxOut_44n[23], nwayMuxOut_45n[23]);
  ND3 I426 (internal_0n[403], nwayMuxOut_46n[23], nwayMuxOut_47n[23], nwayMuxOut_48n[23]);
  NR4 I427 (internal_0n[404], internal_0n[391], internal_0n[392], internal_0n[393], internal_0n[394]);
  NR4 I428 (internal_0n[405], internal_0n[395], internal_0n[396], internal_0n[397], internal_0n[398]);
  NR2 I429 (internal_0n[406], internal_0n[399], internal_0n[400]);
  NR3 I430 (internal_0n[407], internal_0n[401], internal_0n[402], internal_0n[403]);
  ND4 I431 (out_0d[23], internal_0n[404], internal_0n[405], internal_0n[406], internal_0n[407]);
  ND4 I432 (internal_0n[408], nwayMuxOut_0n[24], nwayMuxOut_1n[24], nwayMuxOut_2n[24], nwayMuxOut_3n[24]);
  ND4 I433 (internal_0n[409], nwayMuxOut_4n[24], nwayMuxOut_5n[24], nwayMuxOut_6n[24], nwayMuxOut_7n[24]);
  ND4 I434 (internal_0n[410], nwayMuxOut_8n[24], nwayMuxOut_9n[24], nwayMuxOut_10n[24], nwayMuxOut_11n[24]);
  ND4 I435 (internal_0n[411], nwayMuxOut_12n[24], nwayMuxOut_13n[24], nwayMuxOut_14n[24], nwayMuxOut_15n[24]);
  ND4 I436 (internal_0n[412], nwayMuxOut_16n[24], nwayMuxOut_17n[24], nwayMuxOut_18n[24], nwayMuxOut_19n[24]);
  ND4 I437 (internal_0n[413], nwayMuxOut_20n[24], nwayMuxOut_21n[24], nwayMuxOut_22n[24], nwayMuxOut_23n[24]);
  ND4 I438 (internal_0n[414], nwayMuxOut_24n[24], nwayMuxOut_25n[24], nwayMuxOut_26n[24], nwayMuxOut_27n[24]);
  ND4 I439 (internal_0n[415], nwayMuxOut_28n[24], nwayMuxOut_29n[24], nwayMuxOut_30n[24], nwayMuxOut_31n[24]);
  ND4 I440 (internal_0n[416], nwayMuxOut_32n[24], nwayMuxOut_33n[24], nwayMuxOut_34n[24], nwayMuxOut_35n[24]);
  ND4 I441 (internal_0n[417], nwayMuxOut_36n[24], nwayMuxOut_37n[24], nwayMuxOut_38n[24], nwayMuxOut_39n[24]);
  ND4 I442 (internal_0n[418], nwayMuxOut_40n[24], nwayMuxOut_41n[24], nwayMuxOut_42n[24], nwayMuxOut_43n[24]);
  ND2 I443 (internal_0n[419], nwayMuxOut_44n[24], nwayMuxOut_45n[24]);
  ND3 I444 (internal_0n[420], nwayMuxOut_46n[24], nwayMuxOut_47n[24], nwayMuxOut_48n[24]);
  NR4 I445 (internal_0n[421], internal_0n[408], internal_0n[409], internal_0n[410], internal_0n[411]);
  NR4 I446 (internal_0n[422], internal_0n[412], internal_0n[413], internal_0n[414], internal_0n[415]);
  NR2 I447 (internal_0n[423], internal_0n[416], internal_0n[417]);
  NR3 I448 (internal_0n[424], internal_0n[418], internal_0n[419], internal_0n[420]);
  ND4 I449 (out_0d[24], internal_0n[421], internal_0n[422], internal_0n[423], internal_0n[424]);
  ND4 I450 (internal_0n[425], nwayMuxOut_0n[25], nwayMuxOut_1n[25], nwayMuxOut_2n[25], nwayMuxOut_3n[25]);
  ND4 I451 (internal_0n[426], nwayMuxOut_4n[25], nwayMuxOut_5n[25], nwayMuxOut_6n[25], nwayMuxOut_7n[25]);
  ND4 I452 (internal_0n[427], nwayMuxOut_8n[25], nwayMuxOut_9n[25], nwayMuxOut_10n[25], nwayMuxOut_11n[25]);
  ND4 I453 (internal_0n[428], nwayMuxOut_12n[25], nwayMuxOut_13n[25], nwayMuxOut_14n[25], nwayMuxOut_15n[25]);
  ND4 I454 (internal_0n[429], nwayMuxOut_16n[25], nwayMuxOut_17n[25], nwayMuxOut_18n[25], nwayMuxOut_19n[25]);
  ND4 I455 (internal_0n[430], nwayMuxOut_20n[25], nwayMuxOut_21n[25], nwayMuxOut_22n[25], nwayMuxOut_23n[25]);
  ND4 I456 (internal_0n[431], nwayMuxOut_24n[25], nwayMuxOut_25n[25], nwayMuxOut_26n[25], nwayMuxOut_27n[25]);
  ND4 I457 (internal_0n[432], nwayMuxOut_28n[25], nwayMuxOut_29n[25], nwayMuxOut_30n[25], nwayMuxOut_31n[25]);
  ND4 I458 (internal_0n[433], nwayMuxOut_32n[25], nwayMuxOut_33n[25], nwayMuxOut_34n[25], nwayMuxOut_35n[25]);
  ND4 I459 (internal_0n[434], nwayMuxOut_36n[25], nwayMuxOut_37n[25], nwayMuxOut_38n[25], nwayMuxOut_39n[25]);
  ND4 I460 (internal_0n[435], nwayMuxOut_40n[25], nwayMuxOut_41n[25], nwayMuxOut_42n[25], nwayMuxOut_43n[25]);
  ND2 I461 (internal_0n[436], nwayMuxOut_44n[25], nwayMuxOut_45n[25]);
  ND3 I462 (internal_0n[437], nwayMuxOut_46n[25], nwayMuxOut_47n[25], nwayMuxOut_48n[25]);
  NR4 I463 (internal_0n[438], internal_0n[425], internal_0n[426], internal_0n[427], internal_0n[428]);
  NR4 I464 (internal_0n[439], internal_0n[429], internal_0n[430], internal_0n[431], internal_0n[432]);
  NR2 I465 (internal_0n[440], internal_0n[433], internal_0n[434]);
  NR3 I466 (internal_0n[441], internal_0n[435], internal_0n[436], internal_0n[437]);
  ND4 I467 (out_0d[25], internal_0n[438], internal_0n[439], internal_0n[440], internal_0n[441]);
  ND4 I468 (internal_0n[442], nwayMuxOut_0n[26], nwayMuxOut_1n[26], nwayMuxOut_2n[26], nwayMuxOut_3n[26]);
  ND4 I469 (internal_0n[443], nwayMuxOut_4n[26], nwayMuxOut_5n[26], nwayMuxOut_6n[26], nwayMuxOut_7n[26]);
  ND4 I470 (internal_0n[444], nwayMuxOut_8n[26], nwayMuxOut_9n[26], nwayMuxOut_10n[26], nwayMuxOut_11n[26]);
  ND4 I471 (internal_0n[445], nwayMuxOut_12n[26], nwayMuxOut_13n[26], nwayMuxOut_14n[26], nwayMuxOut_15n[26]);
  ND4 I472 (internal_0n[446], nwayMuxOut_16n[26], nwayMuxOut_17n[26], nwayMuxOut_18n[26], nwayMuxOut_19n[26]);
  ND4 I473 (internal_0n[447], nwayMuxOut_20n[26], nwayMuxOut_21n[26], nwayMuxOut_22n[26], nwayMuxOut_23n[26]);
  ND4 I474 (internal_0n[448], nwayMuxOut_24n[26], nwayMuxOut_25n[26], nwayMuxOut_26n[26], nwayMuxOut_27n[26]);
  ND4 I475 (internal_0n[449], nwayMuxOut_28n[26], nwayMuxOut_29n[26], nwayMuxOut_30n[26], nwayMuxOut_31n[26]);
  ND4 I476 (internal_0n[450], nwayMuxOut_32n[26], nwayMuxOut_33n[26], nwayMuxOut_34n[26], nwayMuxOut_35n[26]);
  ND4 I477 (internal_0n[451], nwayMuxOut_36n[26], nwayMuxOut_37n[26], nwayMuxOut_38n[26], nwayMuxOut_39n[26]);
  ND4 I478 (internal_0n[452], nwayMuxOut_40n[26], nwayMuxOut_41n[26], nwayMuxOut_42n[26], nwayMuxOut_43n[26]);
  ND2 I479 (internal_0n[453], nwayMuxOut_44n[26], nwayMuxOut_45n[26]);
  ND3 I480 (internal_0n[454], nwayMuxOut_46n[26], nwayMuxOut_47n[26], nwayMuxOut_48n[26]);
  NR4 I481 (internal_0n[455], internal_0n[442], internal_0n[443], internal_0n[444], internal_0n[445]);
  NR4 I482 (internal_0n[456], internal_0n[446], internal_0n[447], internal_0n[448], internal_0n[449]);
  NR2 I483 (internal_0n[457], internal_0n[450], internal_0n[451]);
  NR3 I484 (internal_0n[458], internal_0n[452], internal_0n[453], internal_0n[454]);
  ND4 I485 (out_0d[26], internal_0n[455], internal_0n[456], internal_0n[457], internal_0n[458]);
  ND4 I486 (internal_0n[459], nwayMuxOut_0n[27], nwayMuxOut_1n[27], nwayMuxOut_2n[27], nwayMuxOut_3n[27]);
  ND4 I487 (internal_0n[460], nwayMuxOut_4n[27], nwayMuxOut_5n[27], nwayMuxOut_6n[27], nwayMuxOut_7n[27]);
  ND4 I488 (internal_0n[461], nwayMuxOut_8n[27], nwayMuxOut_9n[27], nwayMuxOut_10n[27], nwayMuxOut_11n[27]);
  ND4 I489 (internal_0n[462], nwayMuxOut_12n[27], nwayMuxOut_13n[27], nwayMuxOut_14n[27], nwayMuxOut_15n[27]);
  ND4 I490 (internal_0n[463], nwayMuxOut_16n[27], nwayMuxOut_17n[27], nwayMuxOut_18n[27], nwayMuxOut_19n[27]);
  ND4 I491 (internal_0n[464], nwayMuxOut_20n[27], nwayMuxOut_21n[27], nwayMuxOut_22n[27], nwayMuxOut_23n[27]);
  ND4 I492 (internal_0n[465], nwayMuxOut_24n[27], nwayMuxOut_25n[27], nwayMuxOut_26n[27], nwayMuxOut_27n[27]);
  ND4 I493 (internal_0n[466], nwayMuxOut_28n[27], nwayMuxOut_29n[27], nwayMuxOut_30n[27], nwayMuxOut_31n[27]);
  ND4 I494 (internal_0n[467], nwayMuxOut_32n[27], nwayMuxOut_33n[27], nwayMuxOut_34n[27], nwayMuxOut_35n[27]);
  ND4 I495 (internal_0n[468], nwayMuxOut_36n[27], nwayMuxOut_37n[27], nwayMuxOut_38n[27], nwayMuxOut_39n[27]);
  ND4 I496 (internal_0n[469], nwayMuxOut_40n[27], nwayMuxOut_41n[27], nwayMuxOut_42n[27], nwayMuxOut_43n[27]);
  ND2 I497 (internal_0n[470], nwayMuxOut_44n[27], nwayMuxOut_45n[27]);
  ND3 I498 (internal_0n[471], nwayMuxOut_46n[27], nwayMuxOut_47n[27], nwayMuxOut_48n[27]);
  NR4 I499 (internal_0n[472], internal_0n[459], internal_0n[460], internal_0n[461], internal_0n[462]);
  NR4 I500 (internal_0n[473], internal_0n[463], internal_0n[464], internal_0n[465], internal_0n[466]);
  NR2 I501 (internal_0n[474], internal_0n[467], internal_0n[468]);
  NR3 I502 (internal_0n[475], internal_0n[469], internal_0n[470], internal_0n[471]);
  ND4 I503 (out_0d[27], internal_0n[472], internal_0n[473], internal_0n[474], internal_0n[475]);
  ND4 I504 (internal_0n[476], nwayMuxOut_0n[28], nwayMuxOut_1n[28], nwayMuxOut_2n[28], nwayMuxOut_3n[28]);
  ND4 I505 (internal_0n[477], nwayMuxOut_4n[28], nwayMuxOut_5n[28], nwayMuxOut_6n[28], nwayMuxOut_7n[28]);
  ND4 I506 (internal_0n[478], nwayMuxOut_8n[28], nwayMuxOut_9n[28], nwayMuxOut_10n[28], nwayMuxOut_11n[28]);
  ND4 I507 (internal_0n[479], nwayMuxOut_12n[28], nwayMuxOut_13n[28], nwayMuxOut_14n[28], nwayMuxOut_15n[28]);
  ND4 I508 (internal_0n[480], nwayMuxOut_16n[28], nwayMuxOut_17n[28], nwayMuxOut_18n[28], nwayMuxOut_19n[28]);
  ND4 I509 (internal_0n[481], nwayMuxOut_20n[28], nwayMuxOut_21n[28], nwayMuxOut_22n[28], nwayMuxOut_23n[28]);
  ND4 I510 (internal_0n[482], nwayMuxOut_24n[28], nwayMuxOut_25n[28], nwayMuxOut_26n[28], nwayMuxOut_27n[28]);
  ND4 I511 (internal_0n[483], nwayMuxOut_28n[28], nwayMuxOut_29n[28], nwayMuxOut_30n[28], nwayMuxOut_31n[28]);
  ND4 I512 (internal_0n[484], nwayMuxOut_32n[28], nwayMuxOut_33n[28], nwayMuxOut_34n[28], nwayMuxOut_35n[28]);
  ND4 I513 (internal_0n[485], nwayMuxOut_36n[28], nwayMuxOut_37n[28], nwayMuxOut_38n[28], nwayMuxOut_39n[28]);
  ND4 I514 (internal_0n[486], nwayMuxOut_40n[28], nwayMuxOut_41n[28], nwayMuxOut_42n[28], nwayMuxOut_43n[28]);
  ND2 I515 (internal_0n[487], nwayMuxOut_44n[28], nwayMuxOut_45n[28]);
  ND3 I516 (internal_0n[488], nwayMuxOut_46n[28], nwayMuxOut_47n[28], nwayMuxOut_48n[28]);
  NR4 I517 (internal_0n[489], internal_0n[476], internal_0n[477], internal_0n[478], internal_0n[479]);
  NR4 I518 (internal_0n[490], internal_0n[480], internal_0n[481], internal_0n[482], internal_0n[483]);
  NR2 I519 (internal_0n[491], internal_0n[484], internal_0n[485]);
  NR3 I520 (internal_0n[492], internal_0n[486], internal_0n[487], internal_0n[488]);
  ND4 I521 (out_0d[28], internal_0n[489], internal_0n[490], internal_0n[491], internal_0n[492]);
  ND4 I522 (internal_0n[493], nwayMuxOut_0n[29], nwayMuxOut_1n[29], nwayMuxOut_2n[29], nwayMuxOut_3n[29]);
  ND4 I523 (internal_0n[494], nwayMuxOut_4n[29], nwayMuxOut_5n[29], nwayMuxOut_6n[29], nwayMuxOut_7n[29]);
  ND4 I524 (internal_0n[495], nwayMuxOut_8n[29], nwayMuxOut_9n[29], nwayMuxOut_10n[29], nwayMuxOut_11n[29]);
  ND4 I525 (internal_0n[496], nwayMuxOut_12n[29], nwayMuxOut_13n[29], nwayMuxOut_14n[29], nwayMuxOut_15n[29]);
  ND4 I526 (internal_0n[497], nwayMuxOut_16n[29], nwayMuxOut_17n[29], nwayMuxOut_18n[29], nwayMuxOut_19n[29]);
  ND4 I527 (internal_0n[498], nwayMuxOut_20n[29], nwayMuxOut_21n[29], nwayMuxOut_22n[29], nwayMuxOut_23n[29]);
  ND4 I528 (internal_0n[499], nwayMuxOut_24n[29], nwayMuxOut_25n[29], nwayMuxOut_26n[29], nwayMuxOut_27n[29]);
  ND4 I529 (internal_0n[500], nwayMuxOut_28n[29], nwayMuxOut_29n[29], nwayMuxOut_30n[29], nwayMuxOut_31n[29]);
  ND4 I530 (internal_0n[501], nwayMuxOut_32n[29], nwayMuxOut_33n[29], nwayMuxOut_34n[29], nwayMuxOut_35n[29]);
  ND4 I531 (internal_0n[502], nwayMuxOut_36n[29], nwayMuxOut_37n[29], nwayMuxOut_38n[29], nwayMuxOut_39n[29]);
  ND4 I532 (internal_0n[503], nwayMuxOut_40n[29], nwayMuxOut_41n[29], nwayMuxOut_42n[29], nwayMuxOut_43n[29]);
  ND2 I533 (internal_0n[504], nwayMuxOut_44n[29], nwayMuxOut_45n[29]);
  ND3 I534 (internal_0n[505], nwayMuxOut_46n[29], nwayMuxOut_47n[29], nwayMuxOut_48n[29]);
  NR4 I535 (internal_0n[506], internal_0n[493], internal_0n[494], internal_0n[495], internal_0n[496]);
  NR4 I536 (internal_0n[507], internal_0n[497], internal_0n[498], internal_0n[499], internal_0n[500]);
  NR2 I537 (internal_0n[508], internal_0n[501], internal_0n[502]);
  NR3 I538 (internal_0n[509], internal_0n[503], internal_0n[504], internal_0n[505]);
  ND4 I539 (out_0d[29], internal_0n[506], internal_0n[507], internal_0n[508], internal_0n[509]);
  ND4 I540 (internal_0n[510], nwayMuxOut_0n[30], nwayMuxOut_1n[30], nwayMuxOut_2n[30], nwayMuxOut_3n[30]);
  ND4 I541 (internal_0n[511], nwayMuxOut_4n[30], nwayMuxOut_5n[30], nwayMuxOut_6n[30], nwayMuxOut_7n[30]);
  ND4 I542 (internal_0n[512], nwayMuxOut_8n[30], nwayMuxOut_9n[30], nwayMuxOut_10n[30], nwayMuxOut_11n[30]);
  ND4 I543 (internal_0n[513], nwayMuxOut_12n[30], nwayMuxOut_13n[30], nwayMuxOut_14n[30], nwayMuxOut_15n[30]);
  ND4 I544 (internal_0n[514], nwayMuxOut_16n[30], nwayMuxOut_17n[30], nwayMuxOut_18n[30], nwayMuxOut_19n[30]);
  ND4 I545 (internal_0n[515], nwayMuxOut_20n[30], nwayMuxOut_21n[30], nwayMuxOut_22n[30], nwayMuxOut_23n[30]);
  ND4 I546 (internal_0n[516], nwayMuxOut_24n[30], nwayMuxOut_25n[30], nwayMuxOut_26n[30], nwayMuxOut_27n[30]);
  ND4 I547 (internal_0n[517], nwayMuxOut_28n[30], nwayMuxOut_29n[30], nwayMuxOut_30n[30], nwayMuxOut_31n[30]);
  ND4 I548 (internal_0n[518], nwayMuxOut_32n[30], nwayMuxOut_33n[30], nwayMuxOut_34n[30], nwayMuxOut_35n[30]);
  ND4 I549 (internal_0n[519], nwayMuxOut_36n[30], nwayMuxOut_37n[30], nwayMuxOut_38n[30], nwayMuxOut_39n[30]);
  ND4 I550 (internal_0n[520], nwayMuxOut_40n[30], nwayMuxOut_41n[30], nwayMuxOut_42n[30], nwayMuxOut_43n[30]);
  ND2 I551 (internal_0n[521], nwayMuxOut_44n[30], nwayMuxOut_45n[30]);
  ND3 I552 (internal_0n[522], nwayMuxOut_46n[30], nwayMuxOut_47n[30], nwayMuxOut_48n[30]);
  NR4 I553 (internal_0n[523], internal_0n[510], internal_0n[511], internal_0n[512], internal_0n[513]);
  NR4 I554 (internal_0n[524], internal_0n[514], internal_0n[515], internal_0n[516], internal_0n[517]);
  NR2 I555 (internal_0n[525], internal_0n[518], internal_0n[519]);
  NR3 I556 (internal_0n[526], internal_0n[520], internal_0n[521], internal_0n[522]);
  ND4 I557 (out_0d[30], internal_0n[523], internal_0n[524], internal_0n[525], internal_0n[526]);
  ND4 I558 (internal_0n[527], nwayMuxOut_0n[31], nwayMuxOut_1n[31], nwayMuxOut_2n[31], nwayMuxOut_3n[31]);
  ND4 I559 (internal_0n[528], nwayMuxOut_4n[31], nwayMuxOut_5n[31], nwayMuxOut_6n[31], nwayMuxOut_7n[31]);
  ND4 I560 (internal_0n[529], nwayMuxOut_8n[31], nwayMuxOut_9n[31], nwayMuxOut_10n[31], nwayMuxOut_11n[31]);
  ND4 I561 (internal_0n[530], nwayMuxOut_12n[31], nwayMuxOut_13n[31], nwayMuxOut_14n[31], nwayMuxOut_15n[31]);
  ND4 I562 (internal_0n[531], nwayMuxOut_16n[31], nwayMuxOut_17n[31], nwayMuxOut_18n[31], nwayMuxOut_19n[31]);
  ND4 I563 (internal_0n[532], nwayMuxOut_20n[31], nwayMuxOut_21n[31], nwayMuxOut_22n[31], nwayMuxOut_23n[31]);
  ND4 I564 (internal_0n[533], nwayMuxOut_24n[31], nwayMuxOut_25n[31], nwayMuxOut_26n[31], nwayMuxOut_27n[31]);
  ND4 I565 (internal_0n[534], nwayMuxOut_28n[31], nwayMuxOut_29n[31], nwayMuxOut_30n[31], nwayMuxOut_31n[31]);
  ND4 I566 (internal_0n[535], nwayMuxOut_32n[31], nwayMuxOut_33n[31], nwayMuxOut_34n[31], nwayMuxOut_35n[31]);
  ND4 I567 (internal_0n[536], nwayMuxOut_36n[31], nwayMuxOut_37n[31], nwayMuxOut_38n[31], nwayMuxOut_39n[31]);
  ND4 I568 (internal_0n[537], nwayMuxOut_40n[31], nwayMuxOut_41n[31], nwayMuxOut_42n[31], nwayMuxOut_43n[31]);
  ND2 I569 (internal_0n[538], nwayMuxOut_44n[31], nwayMuxOut_45n[31]);
  ND3 I570 (internal_0n[539], nwayMuxOut_46n[31], nwayMuxOut_47n[31], nwayMuxOut_48n[31]);
  NR4 I571 (internal_0n[540], internal_0n[527], internal_0n[528], internal_0n[529], internal_0n[530]);
  NR4 I572 (internal_0n[541], internal_0n[531], internal_0n[532], internal_0n[533], internal_0n[534]);
  NR2 I573 (internal_0n[542], internal_0n[535], internal_0n[536]);
  NR3 I574 (internal_0n[543], internal_0n[537], internal_0n[538], internal_0n[539]);
  ND4 I575 (out_0d[31], internal_0n[540], internal_0n[541], internal_0n[542], internal_0n[543]);
  ND4 I576 (internal_0n[544], nwayMuxOut_0n[32], nwayMuxOut_1n[32], nwayMuxOut_2n[32], nwayMuxOut_3n[32]);
  ND4 I577 (internal_0n[545], nwayMuxOut_4n[32], nwayMuxOut_5n[32], nwayMuxOut_6n[32], nwayMuxOut_7n[32]);
  ND4 I578 (internal_0n[546], nwayMuxOut_8n[32], nwayMuxOut_9n[32], nwayMuxOut_10n[32], nwayMuxOut_11n[32]);
  ND4 I579 (internal_0n[547], nwayMuxOut_12n[32], nwayMuxOut_13n[32], nwayMuxOut_14n[32], nwayMuxOut_15n[32]);
  ND4 I580 (internal_0n[548], nwayMuxOut_16n[32], nwayMuxOut_17n[32], nwayMuxOut_18n[32], nwayMuxOut_19n[32]);
  ND4 I581 (internal_0n[549], nwayMuxOut_20n[32], nwayMuxOut_21n[32], nwayMuxOut_22n[32], nwayMuxOut_23n[32]);
  ND4 I582 (internal_0n[550], nwayMuxOut_24n[32], nwayMuxOut_25n[32], nwayMuxOut_26n[32], nwayMuxOut_27n[32]);
  ND4 I583 (internal_0n[551], nwayMuxOut_28n[32], nwayMuxOut_29n[32], nwayMuxOut_30n[32], nwayMuxOut_31n[32]);
  ND4 I584 (internal_0n[552], nwayMuxOut_32n[32], nwayMuxOut_33n[32], nwayMuxOut_34n[32], nwayMuxOut_35n[32]);
  ND4 I585 (internal_0n[553], nwayMuxOut_36n[32], nwayMuxOut_37n[32], nwayMuxOut_38n[32], nwayMuxOut_39n[32]);
  ND4 I586 (internal_0n[554], nwayMuxOut_40n[32], nwayMuxOut_41n[32], nwayMuxOut_42n[32], nwayMuxOut_43n[32]);
  ND2 I587 (internal_0n[555], nwayMuxOut_44n[32], nwayMuxOut_45n[32]);
  ND3 I588 (internal_0n[556], nwayMuxOut_46n[32], nwayMuxOut_47n[32], nwayMuxOut_48n[32]);
  NR4 I589 (internal_0n[557], internal_0n[544], internal_0n[545], internal_0n[546], internal_0n[547]);
  NR4 I590 (internal_0n[558], internal_0n[548], internal_0n[549], internal_0n[550], internal_0n[551]);
  NR2 I591 (internal_0n[559], internal_0n[552], internal_0n[553]);
  NR3 I592 (internal_0n[560], internal_0n[554], internal_0n[555], internal_0n[556]);
  ND4 I593 (out_0d[32], internal_0n[557], internal_0n[558], internal_0n[559], internal_0n[560]);
  ND2 I594 (nwayMuxOut_0n[0], inp_0d[0], nwaySelect_0n[0]);
  ND2 I595 (nwayMuxOut_0n[1], inp_0d[1], nwaySelect_0n[0]);
  ND2 I596 (nwayMuxOut_0n[2], inp_0d[2], nwaySelect_0n[0]);
  ND2 I597 (nwayMuxOut_0n[3], inp_0d[3], nwaySelect_0n[0]);
  ND2 I598 (nwayMuxOut_0n[4], inp_0d[4], nwaySelect_0n[0]);
  ND2 I599 (nwayMuxOut_0n[5], inp_0d[5], nwaySelect_0n[0]);
  ND2 I600 (nwayMuxOut_0n[6], inp_0d[6], nwaySelect_0n[0]);
  ND2 I601 (nwayMuxOut_0n[7], inp_0d[7], nwaySelect_0n[0]);
  ND2 I602 (nwayMuxOut_0n[8], inp_0d[8], nwaySelect_0n[0]);
  ND2 I603 (nwayMuxOut_0n[9], inp_0d[9], nwaySelect_0n[0]);
  ND2 I604 (nwayMuxOut_0n[10], inp_0d[10], nwaySelect_0n[0]);
  ND2 I605 (nwayMuxOut_0n[11], inp_0d[11], nwaySelect_0n[0]);
  ND2 I606 (nwayMuxOut_0n[12], inp_0d[12], nwaySelect_0n[0]);
  ND2 I607 (nwayMuxOut_0n[13], inp_0d[13], nwaySelect_0n[0]);
  ND2 I608 (nwayMuxOut_0n[14], inp_0d[14], nwaySelect_0n[0]);
  ND2 I609 (nwayMuxOut_0n[15], inp_0d[15], nwaySelect_0n[0]);
  ND2 I610 (nwayMuxOut_0n[16], inp_0d[16], nwaySelect_0n[0]);
  ND2 I611 (nwayMuxOut_0n[17], inp_0d[17], nwaySelect_0n[0]);
  ND2 I612 (nwayMuxOut_0n[18], inp_0d[18], nwaySelect_0n[0]);
  ND2 I613 (nwayMuxOut_0n[19], inp_0d[19], nwaySelect_0n[0]);
  ND2 I614 (nwayMuxOut_0n[20], inp_0d[20], nwaySelect_0n[0]);
  ND2 I615 (nwayMuxOut_0n[21], inp_0d[21], nwaySelect_0n[0]);
  ND2 I616 (nwayMuxOut_0n[22], inp_0d[22], nwaySelect_0n[0]);
  ND2 I617 (nwayMuxOut_0n[23], inp_0d[23], nwaySelect_0n[0]);
  ND2 I618 (nwayMuxOut_0n[24], inp_0d[24], nwaySelect_0n[0]);
  ND2 I619 (nwayMuxOut_0n[25], inp_0d[25], nwaySelect_0n[0]);
  ND2 I620 (nwayMuxOut_0n[26], inp_0d[26], nwaySelect_0n[0]);
  ND2 I621 (nwayMuxOut_0n[27], inp_0d[27], nwaySelect_0n[0]);
  ND2 I622 (nwayMuxOut_0n[28], inp_0d[28], nwaySelect_0n[0]);
  ND2 I623 (nwayMuxOut_0n[29], inp_0d[29], nwaySelect_0n[0]);
  ND2 I624 (nwayMuxOut_0n[30], inp_0d[30], nwaySelect_0n[0]);
  ND2 I625 (nwayMuxOut_0n[31], inp_0d[31], nwaySelect_0n[0]);
  ND2 I626 (nwayMuxOut_0n[32], inp_0d[32], nwaySelect_0n[0]);
  ND2 I627 (nwayMuxOut_1n[0], inp_1d[0], nwaySelect_0n[1]);
  ND2 I628 (nwayMuxOut_1n[1], inp_1d[1], nwaySelect_0n[1]);
  ND2 I629 (nwayMuxOut_1n[2], inp_1d[2], nwaySelect_0n[1]);
  ND2 I630 (nwayMuxOut_1n[3], inp_1d[3], nwaySelect_0n[1]);
  ND2 I631 (nwayMuxOut_1n[4], inp_1d[4], nwaySelect_0n[1]);
  ND2 I632 (nwayMuxOut_1n[5], inp_1d[5], nwaySelect_0n[1]);
  ND2 I633 (nwayMuxOut_1n[6], inp_1d[6], nwaySelect_0n[1]);
  ND2 I634 (nwayMuxOut_1n[7], inp_1d[7], nwaySelect_0n[1]);
  ND2 I635 (nwayMuxOut_1n[8], inp_1d[8], nwaySelect_0n[1]);
  ND2 I636 (nwayMuxOut_1n[9], inp_1d[9], nwaySelect_0n[1]);
  ND2 I637 (nwayMuxOut_1n[10], inp_1d[10], nwaySelect_0n[1]);
  ND2 I638 (nwayMuxOut_1n[11], inp_1d[11], nwaySelect_0n[1]);
  ND2 I639 (nwayMuxOut_1n[12], inp_1d[12], nwaySelect_0n[1]);
  ND2 I640 (nwayMuxOut_1n[13], inp_1d[13], nwaySelect_0n[1]);
  ND2 I641 (nwayMuxOut_1n[14], inp_1d[14], nwaySelect_0n[1]);
  ND2 I642 (nwayMuxOut_1n[15], inp_1d[15], nwaySelect_0n[1]);
  ND2 I643 (nwayMuxOut_1n[16], inp_1d[16], nwaySelect_0n[1]);
  ND2 I644 (nwayMuxOut_1n[17], inp_1d[17], nwaySelect_0n[1]);
  ND2 I645 (nwayMuxOut_1n[18], inp_1d[18], nwaySelect_0n[1]);
  ND2 I646 (nwayMuxOut_1n[19], inp_1d[19], nwaySelect_0n[1]);
  ND2 I647 (nwayMuxOut_1n[20], inp_1d[20], nwaySelect_0n[1]);
  ND2 I648 (nwayMuxOut_1n[21], inp_1d[21], nwaySelect_0n[1]);
  ND2 I649 (nwayMuxOut_1n[22], inp_1d[22], nwaySelect_0n[1]);
  ND2 I650 (nwayMuxOut_1n[23], inp_1d[23], nwaySelect_0n[1]);
  ND2 I651 (nwayMuxOut_1n[24], inp_1d[24], nwaySelect_0n[1]);
  ND2 I652 (nwayMuxOut_1n[25], inp_1d[25], nwaySelect_0n[1]);
  ND2 I653 (nwayMuxOut_1n[26], inp_1d[26], nwaySelect_0n[1]);
  ND2 I654 (nwayMuxOut_1n[27], inp_1d[27], nwaySelect_0n[1]);
  ND2 I655 (nwayMuxOut_1n[28], inp_1d[28], nwaySelect_0n[1]);
  ND2 I656 (nwayMuxOut_1n[29], inp_1d[29], nwaySelect_0n[1]);
  ND2 I657 (nwayMuxOut_1n[30], inp_1d[30], nwaySelect_0n[1]);
  ND2 I658 (nwayMuxOut_1n[31], inp_1d[31], nwaySelect_0n[1]);
  ND2 I659 (nwayMuxOut_1n[32], inp_1d[32], nwaySelect_0n[1]);
  ND2 I660 (nwayMuxOut_2n[0], inp_2d[0], nwaySelect_0n[2]);
  ND2 I661 (nwayMuxOut_2n[1], inp_2d[1], nwaySelect_0n[2]);
  ND2 I662 (nwayMuxOut_2n[2], inp_2d[2], nwaySelect_0n[2]);
  ND2 I663 (nwayMuxOut_2n[3], inp_2d[3], nwaySelect_0n[2]);
  ND2 I664 (nwayMuxOut_2n[4], inp_2d[4], nwaySelect_0n[2]);
  ND2 I665 (nwayMuxOut_2n[5], inp_2d[5], nwaySelect_0n[2]);
  ND2 I666 (nwayMuxOut_2n[6], inp_2d[6], nwaySelect_0n[2]);
  ND2 I667 (nwayMuxOut_2n[7], inp_2d[7], nwaySelect_0n[2]);
  ND2 I668 (nwayMuxOut_2n[8], inp_2d[8], nwaySelect_0n[2]);
  ND2 I669 (nwayMuxOut_2n[9], inp_2d[9], nwaySelect_0n[2]);
  ND2 I670 (nwayMuxOut_2n[10], inp_2d[10], nwaySelect_0n[2]);
  ND2 I671 (nwayMuxOut_2n[11], inp_2d[11], nwaySelect_0n[2]);
  ND2 I672 (nwayMuxOut_2n[12], inp_2d[12], nwaySelect_0n[2]);
  ND2 I673 (nwayMuxOut_2n[13], inp_2d[13], nwaySelect_0n[2]);
  ND2 I674 (nwayMuxOut_2n[14], inp_2d[14], nwaySelect_0n[2]);
  ND2 I675 (nwayMuxOut_2n[15], inp_2d[15], nwaySelect_0n[2]);
  ND2 I676 (nwayMuxOut_2n[16], inp_2d[16], nwaySelect_0n[2]);
  ND2 I677 (nwayMuxOut_2n[17], inp_2d[17], nwaySelect_0n[2]);
  ND2 I678 (nwayMuxOut_2n[18], inp_2d[18], nwaySelect_0n[2]);
  ND2 I679 (nwayMuxOut_2n[19], inp_2d[19], nwaySelect_0n[2]);
  ND2 I680 (nwayMuxOut_2n[20], inp_2d[20], nwaySelect_0n[2]);
  ND2 I681 (nwayMuxOut_2n[21], inp_2d[21], nwaySelect_0n[2]);
  ND2 I682 (nwayMuxOut_2n[22], inp_2d[22], nwaySelect_0n[2]);
  ND2 I683 (nwayMuxOut_2n[23], inp_2d[23], nwaySelect_0n[2]);
  ND2 I684 (nwayMuxOut_2n[24], inp_2d[24], nwaySelect_0n[2]);
  ND2 I685 (nwayMuxOut_2n[25], inp_2d[25], nwaySelect_0n[2]);
  ND2 I686 (nwayMuxOut_2n[26], inp_2d[26], nwaySelect_0n[2]);
  ND2 I687 (nwayMuxOut_2n[27], inp_2d[27], nwaySelect_0n[2]);
  ND2 I688 (nwayMuxOut_2n[28], inp_2d[28], nwaySelect_0n[2]);
  ND2 I689 (nwayMuxOut_2n[29], inp_2d[29], nwaySelect_0n[2]);
  ND2 I690 (nwayMuxOut_2n[30], inp_2d[30], nwaySelect_0n[2]);
  ND2 I691 (nwayMuxOut_2n[31], inp_2d[31], nwaySelect_0n[2]);
  ND2 I692 (nwayMuxOut_2n[32], inp_2d[32], nwaySelect_0n[2]);
  ND2 I693 (nwayMuxOut_3n[0], inp_3d[0], nwaySelect_0n[3]);
  ND2 I694 (nwayMuxOut_3n[1], inp_3d[1], nwaySelect_0n[3]);
  ND2 I695 (nwayMuxOut_3n[2], inp_3d[2], nwaySelect_0n[3]);
  ND2 I696 (nwayMuxOut_3n[3], inp_3d[3], nwaySelect_0n[3]);
  ND2 I697 (nwayMuxOut_3n[4], inp_3d[4], nwaySelect_0n[3]);
  ND2 I698 (nwayMuxOut_3n[5], inp_3d[5], nwaySelect_0n[3]);
  ND2 I699 (nwayMuxOut_3n[6], inp_3d[6], nwaySelect_0n[3]);
  ND2 I700 (nwayMuxOut_3n[7], inp_3d[7], nwaySelect_0n[3]);
  ND2 I701 (nwayMuxOut_3n[8], inp_3d[8], nwaySelect_0n[3]);
  ND2 I702 (nwayMuxOut_3n[9], inp_3d[9], nwaySelect_0n[3]);
  ND2 I703 (nwayMuxOut_3n[10], inp_3d[10], nwaySelect_0n[3]);
  ND2 I704 (nwayMuxOut_3n[11], inp_3d[11], nwaySelect_0n[3]);
  ND2 I705 (nwayMuxOut_3n[12], inp_3d[12], nwaySelect_0n[3]);
  ND2 I706 (nwayMuxOut_3n[13], inp_3d[13], nwaySelect_0n[3]);
  ND2 I707 (nwayMuxOut_3n[14], inp_3d[14], nwaySelect_0n[3]);
  ND2 I708 (nwayMuxOut_3n[15], inp_3d[15], nwaySelect_0n[3]);
  ND2 I709 (nwayMuxOut_3n[16], inp_3d[16], nwaySelect_0n[3]);
  ND2 I710 (nwayMuxOut_3n[17], inp_3d[17], nwaySelect_0n[3]);
  ND2 I711 (nwayMuxOut_3n[18], inp_3d[18], nwaySelect_0n[3]);
  ND2 I712 (nwayMuxOut_3n[19], inp_3d[19], nwaySelect_0n[3]);
  ND2 I713 (nwayMuxOut_3n[20], inp_3d[20], nwaySelect_0n[3]);
  ND2 I714 (nwayMuxOut_3n[21], inp_3d[21], nwaySelect_0n[3]);
  ND2 I715 (nwayMuxOut_3n[22], inp_3d[22], nwaySelect_0n[3]);
  ND2 I716 (nwayMuxOut_3n[23], inp_3d[23], nwaySelect_0n[3]);
  ND2 I717 (nwayMuxOut_3n[24], inp_3d[24], nwaySelect_0n[3]);
  ND2 I718 (nwayMuxOut_3n[25], inp_3d[25], nwaySelect_0n[3]);
  ND2 I719 (nwayMuxOut_3n[26], inp_3d[26], nwaySelect_0n[3]);
  ND2 I720 (nwayMuxOut_3n[27], inp_3d[27], nwaySelect_0n[3]);
  ND2 I721 (nwayMuxOut_3n[28], inp_3d[28], nwaySelect_0n[3]);
  ND2 I722 (nwayMuxOut_3n[29], inp_3d[29], nwaySelect_0n[3]);
  ND2 I723 (nwayMuxOut_3n[30], inp_3d[30], nwaySelect_0n[3]);
  ND2 I724 (nwayMuxOut_3n[31], inp_3d[31], nwaySelect_0n[3]);
  ND2 I725 (nwayMuxOut_3n[32], inp_3d[32], nwaySelect_0n[3]);
  ND2 I726 (nwayMuxOut_4n[0], inp_4d[0], nwaySelect_0n[4]);
  ND2 I727 (nwayMuxOut_4n[1], inp_4d[1], nwaySelect_0n[4]);
  ND2 I728 (nwayMuxOut_4n[2], inp_4d[2], nwaySelect_0n[4]);
  ND2 I729 (nwayMuxOut_4n[3], inp_4d[3], nwaySelect_0n[4]);
  ND2 I730 (nwayMuxOut_4n[4], inp_4d[4], nwaySelect_0n[4]);
  ND2 I731 (nwayMuxOut_4n[5], inp_4d[5], nwaySelect_0n[4]);
  ND2 I732 (nwayMuxOut_4n[6], inp_4d[6], nwaySelect_0n[4]);
  ND2 I733 (nwayMuxOut_4n[7], inp_4d[7], nwaySelect_0n[4]);
  ND2 I734 (nwayMuxOut_4n[8], inp_4d[8], nwaySelect_0n[4]);
  ND2 I735 (nwayMuxOut_4n[9], inp_4d[9], nwaySelect_0n[4]);
  ND2 I736 (nwayMuxOut_4n[10], inp_4d[10], nwaySelect_0n[4]);
  ND2 I737 (nwayMuxOut_4n[11], inp_4d[11], nwaySelect_0n[4]);
  ND2 I738 (nwayMuxOut_4n[12], inp_4d[12], nwaySelect_0n[4]);
  ND2 I739 (nwayMuxOut_4n[13], inp_4d[13], nwaySelect_0n[4]);
  ND2 I740 (nwayMuxOut_4n[14], inp_4d[14], nwaySelect_0n[4]);
  ND2 I741 (nwayMuxOut_4n[15], inp_4d[15], nwaySelect_0n[4]);
  ND2 I742 (nwayMuxOut_4n[16], inp_4d[16], nwaySelect_0n[4]);
  ND2 I743 (nwayMuxOut_4n[17], inp_4d[17], nwaySelect_0n[4]);
  ND2 I744 (nwayMuxOut_4n[18], inp_4d[18], nwaySelect_0n[4]);
  ND2 I745 (nwayMuxOut_4n[19], inp_4d[19], nwaySelect_0n[4]);
  ND2 I746 (nwayMuxOut_4n[20], inp_4d[20], nwaySelect_0n[4]);
  ND2 I747 (nwayMuxOut_4n[21], inp_4d[21], nwaySelect_0n[4]);
  ND2 I748 (nwayMuxOut_4n[22], inp_4d[22], nwaySelect_0n[4]);
  ND2 I749 (nwayMuxOut_4n[23], inp_4d[23], nwaySelect_0n[4]);
  ND2 I750 (nwayMuxOut_4n[24], inp_4d[24], nwaySelect_0n[4]);
  ND2 I751 (nwayMuxOut_4n[25], inp_4d[25], nwaySelect_0n[4]);
  ND2 I752 (nwayMuxOut_4n[26], inp_4d[26], nwaySelect_0n[4]);
  ND2 I753 (nwayMuxOut_4n[27], inp_4d[27], nwaySelect_0n[4]);
  ND2 I754 (nwayMuxOut_4n[28], inp_4d[28], nwaySelect_0n[4]);
  ND2 I755 (nwayMuxOut_4n[29], inp_4d[29], nwaySelect_0n[4]);
  ND2 I756 (nwayMuxOut_4n[30], inp_4d[30], nwaySelect_0n[4]);
  ND2 I757 (nwayMuxOut_4n[31], inp_4d[31], nwaySelect_0n[4]);
  ND2 I758 (nwayMuxOut_4n[32], inp_4d[32], nwaySelect_0n[4]);
  ND2 I759 (nwayMuxOut_5n[0], inp_5d[0], nwaySelect_0n[5]);
  ND2 I760 (nwayMuxOut_5n[1], inp_5d[1], nwaySelect_0n[5]);
  ND2 I761 (nwayMuxOut_5n[2], inp_5d[2], nwaySelect_0n[5]);
  ND2 I762 (nwayMuxOut_5n[3], inp_5d[3], nwaySelect_0n[5]);
  ND2 I763 (nwayMuxOut_5n[4], inp_5d[4], nwaySelect_0n[5]);
  ND2 I764 (nwayMuxOut_5n[5], inp_5d[5], nwaySelect_0n[5]);
  ND2 I765 (nwayMuxOut_5n[6], inp_5d[6], nwaySelect_0n[5]);
  ND2 I766 (nwayMuxOut_5n[7], inp_5d[7], nwaySelect_0n[5]);
  ND2 I767 (nwayMuxOut_5n[8], inp_5d[8], nwaySelect_0n[5]);
  ND2 I768 (nwayMuxOut_5n[9], inp_5d[9], nwaySelect_0n[5]);
  ND2 I769 (nwayMuxOut_5n[10], inp_5d[10], nwaySelect_0n[5]);
  ND2 I770 (nwayMuxOut_5n[11], inp_5d[11], nwaySelect_0n[5]);
  ND2 I771 (nwayMuxOut_5n[12], inp_5d[12], nwaySelect_0n[5]);
  ND2 I772 (nwayMuxOut_5n[13], inp_5d[13], nwaySelect_0n[5]);
  ND2 I773 (nwayMuxOut_5n[14], inp_5d[14], nwaySelect_0n[5]);
  ND2 I774 (nwayMuxOut_5n[15], inp_5d[15], nwaySelect_0n[5]);
  ND2 I775 (nwayMuxOut_5n[16], inp_5d[16], nwaySelect_0n[5]);
  ND2 I776 (nwayMuxOut_5n[17], inp_5d[17], nwaySelect_0n[5]);
  ND2 I777 (nwayMuxOut_5n[18], inp_5d[18], nwaySelect_0n[5]);
  ND2 I778 (nwayMuxOut_5n[19], inp_5d[19], nwaySelect_0n[5]);
  ND2 I779 (nwayMuxOut_5n[20], inp_5d[20], nwaySelect_0n[5]);
  ND2 I780 (nwayMuxOut_5n[21], inp_5d[21], nwaySelect_0n[5]);
  ND2 I781 (nwayMuxOut_5n[22], inp_5d[22], nwaySelect_0n[5]);
  ND2 I782 (nwayMuxOut_5n[23], inp_5d[23], nwaySelect_0n[5]);
  ND2 I783 (nwayMuxOut_5n[24], inp_5d[24], nwaySelect_0n[5]);
  ND2 I784 (nwayMuxOut_5n[25], inp_5d[25], nwaySelect_0n[5]);
  ND2 I785 (nwayMuxOut_5n[26], inp_5d[26], nwaySelect_0n[5]);
  ND2 I786 (nwayMuxOut_5n[27], inp_5d[27], nwaySelect_0n[5]);
  ND2 I787 (nwayMuxOut_5n[28], inp_5d[28], nwaySelect_0n[5]);
  ND2 I788 (nwayMuxOut_5n[29], inp_5d[29], nwaySelect_0n[5]);
  ND2 I789 (nwayMuxOut_5n[30], inp_5d[30], nwaySelect_0n[5]);
  ND2 I790 (nwayMuxOut_5n[31], inp_5d[31], nwaySelect_0n[5]);
  ND2 I791 (nwayMuxOut_5n[32], inp_5d[32], nwaySelect_0n[5]);
  ND2 I792 (nwayMuxOut_6n[0], inp_6d[0], nwaySelect_0n[6]);
  ND2 I793 (nwayMuxOut_6n[1], inp_6d[1], nwaySelect_0n[6]);
  ND2 I794 (nwayMuxOut_6n[2], inp_6d[2], nwaySelect_0n[6]);
  ND2 I795 (nwayMuxOut_6n[3], inp_6d[3], nwaySelect_0n[6]);
  ND2 I796 (nwayMuxOut_6n[4], inp_6d[4], nwaySelect_0n[6]);
  ND2 I797 (nwayMuxOut_6n[5], inp_6d[5], nwaySelect_0n[6]);
  ND2 I798 (nwayMuxOut_6n[6], inp_6d[6], nwaySelect_0n[6]);
  ND2 I799 (nwayMuxOut_6n[7], inp_6d[7], nwaySelect_0n[6]);
  ND2 I800 (nwayMuxOut_6n[8], inp_6d[8], nwaySelect_0n[6]);
  ND2 I801 (nwayMuxOut_6n[9], inp_6d[9], nwaySelect_0n[6]);
  ND2 I802 (nwayMuxOut_6n[10], inp_6d[10], nwaySelect_0n[6]);
  ND2 I803 (nwayMuxOut_6n[11], inp_6d[11], nwaySelect_0n[6]);
  ND2 I804 (nwayMuxOut_6n[12], inp_6d[12], nwaySelect_0n[6]);
  ND2 I805 (nwayMuxOut_6n[13], inp_6d[13], nwaySelect_0n[6]);
  ND2 I806 (nwayMuxOut_6n[14], inp_6d[14], nwaySelect_0n[6]);
  ND2 I807 (nwayMuxOut_6n[15], inp_6d[15], nwaySelect_0n[6]);
  ND2 I808 (nwayMuxOut_6n[16], inp_6d[16], nwaySelect_0n[6]);
  ND2 I809 (nwayMuxOut_6n[17], inp_6d[17], nwaySelect_0n[6]);
  ND2 I810 (nwayMuxOut_6n[18], inp_6d[18], nwaySelect_0n[6]);
  ND2 I811 (nwayMuxOut_6n[19], inp_6d[19], nwaySelect_0n[6]);
  ND2 I812 (nwayMuxOut_6n[20], inp_6d[20], nwaySelect_0n[6]);
  ND2 I813 (nwayMuxOut_6n[21], inp_6d[21], nwaySelect_0n[6]);
  ND2 I814 (nwayMuxOut_6n[22], inp_6d[22], nwaySelect_0n[6]);
  ND2 I815 (nwayMuxOut_6n[23], inp_6d[23], nwaySelect_0n[6]);
  ND2 I816 (nwayMuxOut_6n[24], inp_6d[24], nwaySelect_0n[6]);
  ND2 I817 (nwayMuxOut_6n[25], inp_6d[25], nwaySelect_0n[6]);
  ND2 I818 (nwayMuxOut_6n[26], inp_6d[26], nwaySelect_0n[6]);
  ND2 I819 (nwayMuxOut_6n[27], inp_6d[27], nwaySelect_0n[6]);
  ND2 I820 (nwayMuxOut_6n[28], inp_6d[28], nwaySelect_0n[6]);
  ND2 I821 (nwayMuxOut_6n[29], inp_6d[29], nwaySelect_0n[6]);
  ND2 I822 (nwayMuxOut_6n[30], inp_6d[30], nwaySelect_0n[6]);
  ND2 I823 (nwayMuxOut_6n[31], inp_6d[31], nwaySelect_0n[6]);
  ND2 I824 (nwayMuxOut_6n[32], inp_6d[32], nwaySelect_0n[6]);
  ND2 I825 (nwayMuxOut_7n[0], inp_7d[0], nwaySelect_0n[7]);
  ND2 I826 (nwayMuxOut_7n[1], inp_7d[1], nwaySelect_0n[7]);
  ND2 I827 (nwayMuxOut_7n[2], inp_7d[2], nwaySelect_0n[7]);
  ND2 I828 (nwayMuxOut_7n[3], inp_7d[3], nwaySelect_0n[7]);
  ND2 I829 (nwayMuxOut_7n[4], inp_7d[4], nwaySelect_0n[7]);
  ND2 I830 (nwayMuxOut_7n[5], inp_7d[5], nwaySelect_0n[7]);
  ND2 I831 (nwayMuxOut_7n[6], inp_7d[6], nwaySelect_0n[7]);
  ND2 I832 (nwayMuxOut_7n[7], inp_7d[7], nwaySelect_0n[7]);
  ND2 I833 (nwayMuxOut_7n[8], inp_7d[8], nwaySelect_0n[7]);
  ND2 I834 (nwayMuxOut_7n[9], inp_7d[9], nwaySelect_0n[7]);
  ND2 I835 (nwayMuxOut_7n[10], inp_7d[10], nwaySelect_0n[7]);
  ND2 I836 (nwayMuxOut_7n[11], inp_7d[11], nwaySelect_0n[7]);
  ND2 I837 (nwayMuxOut_7n[12], inp_7d[12], nwaySelect_0n[7]);
  ND2 I838 (nwayMuxOut_7n[13], inp_7d[13], nwaySelect_0n[7]);
  ND2 I839 (nwayMuxOut_7n[14], inp_7d[14], nwaySelect_0n[7]);
  ND2 I840 (nwayMuxOut_7n[15], inp_7d[15], nwaySelect_0n[7]);
  ND2 I841 (nwayMuxOut_7n[16], inp_7d[16], nwaySelect_0n[7]);
  ND2 I842 (nwayMuxOut_7n[17], inp_7d[17], nwaySelect_0n[7]);
  ND2 I843 (nwayMuxOut_7n[18], inp_7d[18], nwaySelect_0n[7]);
  ND2 I844 (nwayMuxOut_7n[19], inp_7d[19], nwaySelect_0n[7]);
  ND2 I845 (nwayMuxOut_7n[20], inp_7d[20], nwaySelect_0n[7]);
  ND2 I846 (nwayMuxOut_7n[21], inp_7d[21], nwaySelect_0n[7]);
  ND2 I847 (nwayMuxOut_7n[22], inp_7d[22], nwaySelect_0n[7]);
  ND2 I848 (nwayMuxOut_7n[23], inp_7d[23], nwaySelect_0n[7]);
  ND2 I849 (nwayMuxOut_7n[24], inp_7d[24], nwaySelect_0n[7]);
  ND2 I850 (nwayMuxOut_7n[25], inp_7d[25], nwaySelect_0n[7]);
  ND2 I851 (nwayMuxOut_7n[26], inp_7d[26], nwaySelect_0n[7]);
  ND2 I852 (nwayMuxOut_7n[27], inp_7d[27], nwaySelect_0n[7]);
  ND2 I853 (nwayMuxOut_7n[28], inp_7d[28], nwaySelect_0n[7]);
  ND2 I854 (nwayMuxOut_7n[29], inp_7d[29], nwaySelect_0n[7]);
  ND2 I855 (nwayMuxOut_7n[30], inp_7d[30], nwaySelect_0n[7]);
  ND2 I856 (nwayMuxOut_7n[31], inp_7d[31], nwaySelect_0n[7]);
  ND2 I857 (nwayMuxOut_7n[32], inp_7d[32], nwaySelect_0n[7]);
  ND2 I858 (nwayMuxOut_8n[0], inp_8d[0], nwaySelect_0n[8]);
  ND2 I859 (nwayMuxOut_8n[1], inp_8d[1], nwaySelect_0n[8]);
  ND2 I860 (nwayMuxOut_8n[2], inp_8d[2], nwaySelect_0n[8]);
  ND2 I861 (nwayMuxOut_8n[3], inp_8d[3], nwaySelect_0n[8]);
  ND2 I862 (nwayMuxOut_8n[4], inp_8d[4], nwaySelect_0n[8]);
  ND2 I863 (nwayMuxOut_8n[5], inp_8d[5], nwaySelect_0n[8]);
  ND2 I864 (nwayMuxOut_8n[6], inp_8d[6], nwaySelect_0n[8]);
  ND2 I865 (nwayMuxOut_8n[7], inp_8d[7], nwaySelect_0n[8]);
  ND2 I866 (nwayMuxOut_8n[8], inp_8d[8], nwaySelect_0n[8]);
  ND2 I867 (nwayMuxOut_8n[9], inp_8d[9], nwaySelect_0n[8]);
  ND2 I868 (nwayMuxOut_8n[10], inp_8d[10], nwaySelect_0n[8]);
  ND2 I869 (nwayMuxOut_8n[11], inp_8d[11], nwaySelect_0n[8]);
  ND2 I870 (nwayMuxOut_8n[12], inp_8d[12], nwaySelect_0n[8]);
  ND2 I871 (nwayMuxOut_8n[13], inp_8d[13], nwaySelect_0n[8]);
  ND2 I872 (nwayMuxOut_8n[14], inp_8d[14], nwaySelect_0n[8]);
  ND2 I873 (nwayMuxOut_8n[15], inp_8d[15], nwaySelect_0n[8]);
  ND2 I874 (nwayMuxOut_8n[16], inp_8d[16], nwaySelect_0n[8]);
  ND2 I875 (nwayMuxOut_8n[17], inp_8d[17], nwaySelect_0n[8]);
  ND2 I876 (nwayMuxOut_8n[18], inp_8d[18], nwaySelect_0n[8]);
  ND2 I877 (nwayMuxOut_8n[19], inp_8d[19], nwaySelect_0n[8]);
  ND2 I878 (nwayMuxOut_8n[20], inp_8d[20], nwaySelect_0n[8]);
  ND2 I879 (nwayMuxOut_8n[21], inp_8d[21], nwaySelect_0n[8]);
  ND2 I880 (nwayMuxOut_8n[22], inp_8d[22], nwaySelect_0n[8]);
  ND2 I881 (nwayMuxOut_8n[23], inp_8d[23], nwaySelect_0n[8]);
  ND2 I882 (nwayMuxOut_8n[24], inp_8d[24], nwaySelect_0n[8]);
  ND2 I883 (nwayMuxOut_8n[25], inp_8d[25], nwaySelect_0n[8]);
  ND2 I884 (nwayMuxOut_8n[26], inp_8d[26], nwaySelect_0n[8]);
  ND2 I885 (nwayMuxOut_8n[27], inp_8d[27], nwaySelect_0n[8]);
  ND2 I886 (nwayMuxOut_8n[28], inp_8d[28], nwaySelect_0n[8]);
  ND2 I887 (nwayMuxOut_8n[29], inp_8d[29], nwaySelect_0n[8]);
  ND2 I888 (nwayMuxOut_8n[30], inp_8d[30], nwaySelect_0n[8]);
  ND2 I889 (nwayMuxOut_8n[31], inp_8d[31], nwaySelect_0n[8]);
  ND2 I890 (nwayMuxOut_8n[32], inp_8d[32], nwaySelect_0n[8]);
  ND2 I891 (nwayMuxOut_9n[0], inp_9d[0], nwaySelect_0n[9]);
  ND2 I892 (nwayMuxOut_9n[1], inp_9d[1], nwaySelect_0n[9]);
  ND2 I893 (nwayMuxOut_9n[2], inp_9d[2], nwaySelect_0n[9]);
  ND2 I894 (nwayMuxOut_9n[3], inp_9d[3], nwaySelect_0n[9]);
  ND2 I895 (nwayMuxOut_9n[4], inp_9d[4], nwaySelect_0n[9]);
  ND2 I896 (nwayMuxOut_9n[5], inp_9d[5], nwaySelect_0n[9]);
  ND2 I897 (nwayMuxOut_9n[6], inp_9d[6], nwaySelect_0n[9]);
  ND2 I898 (nwayMuxOut_9n[7], inp_9d[7], nwaySelect_0n[9]);
  ND2 I899 (nwayMuxOut_9n[8], inp_9d[8], nwaySelect_0n[9]);
  ND2 I900 (nwayMuxOut_9n[9], inp_9d[9], nwaySelect_0n[9]);
  ND2 I901 (nwayMuxOut_9n[10], inp_9d[10], nwaySelect_0n[9]);
  ND2 I902 (nwayMuxOut_9n[11], inp_9d[11], nwaySelect_0n[9]);
  ND2 I903 (nwayMuxOut_9n[12], inp_9d[12], nwaySelect_0n[9]);
  ND2 I904 (nwayMuxOut_9n[13], inp_9d[13], nwaySelect_0n[9]);
  ND2 I905 (nwayMuxOut_9n[14], inp_9d[14], nwaySelect_0n[9]);
  ND2 I906 (nwayMuxOut_9n[15], inp_9d[15], nwaySelect_0n[9]);
  ND2 I907 (nwayMuxOut_9n[16], inp_9d[16], nwaySelect_0n[9]);
  ND2 I908 (nwayMuxOut_9n[17], inp_9d[17], nwaySelect_0n[9]);
  ND2 I909 (nwayMuxOut_9n[18], inp_9d[18], nwaySelect_0n[9]);
  ND2 I910 (nwayMuxOut_9n[19], inp_9d[19], nwaySelect_0n[9]);
  ND2 I911 (nwayMuxOut_9n[20], inp_9d[20], nwaySelect_0n[9]);
  ND2 I912 (nwayMuxOut_9n[21], inp_9d[21], nwaySelect_0n[9]);
  ND2 I913 (nwayMuxOut_9n[22], inp_9d[22], nwaySelect_0n[9]);
  ND2 I914 (nwayMuxOut_9n[23], inp_9d[23], nwaySelect_0n[9]);
  ND2 I915 (nwayMuxOut_9n[24], inp_9d[24], nwaySelect_0n[9]);
  ND2 I916 (nwayMuxOut_9n[25], inp_9d[25], nwaySelect_0n[9]);
  ND2 I917 (nwayMuxOut_9n[26], inp_9d[26], nwaySelect_0n[9]);
  ND2 I918 (nwayMuxOut_9n[27], inp_9d[27], nwaySelect_0n[9]);
  ND2 I919 (nwayMuxOut_9n[28], inp_9d[28], nwaySelect_0n[9]);
  ND2 I920 (nwayMuxOut_9n[29], inp_9d[29], nwaySelect_0n[9]);
  ND2 I921 (nwayMuxOut_9n[30], inp_9d[30], nwaySelect_0n[9]);
  ND2 I922 (nwayMuxOut_9n[31], inp_9d[31], nwaySelect_0n[9]);
  ND2 I923 (nwayMuxOut_9n[32], inp_9d[32], nwaySelect_0n[9]);
  ND2 I924 (nwayMuxOut_10n[0], inp_10d[0], nwaySelect_0n[10]);
  ND2 I925 (nwayMuxOut_10n[1], inp_10d[1], nwaySelect_0n[10]);
  ND2 I926 (nwayMuxOut_10n[2], inp_10d[2], nwaySelect_0n[10]);
  ND2 I927 (nwayMuxOut_10n[3], inp_10d[3], nwaySelect_0n[10]);
  ND2 I928 (nwayMuxOut_10n[4], inp_10d[4], nwaySelect_0n[10]);
  ND2 I929 (nwayMuxOut_10n[5], inp_10d[5], nwaySelect_0n[10]);
  ND2 I930 (nwayMuxOut_10n[6], inp_10d[6], nwaySelect_0n[10]);
  ND2 I931 (nwayMuxOut_10n[7], inp_10d[7], nwaySelect_0n[10]);
  ND2 I932 (nwayMuxOut_10n[8], inp_10d[8], nwaySelect_0n[10]);
  ND2 I933 (nwayMuxOut_10n[9], inp_10d[9], nwaySelect_0n[10]);
  ND2 I934 (nwayMuxOut_10n[10], inp_10d[10], nwaySelect_0n[10]);
  ND2 I935 (nwayMuxOut_10n[11], inp_10d[11], nwaySelect_0n[10]);
  ND2 I936 (nwayMuxOut_10n[12], inp_10d[12], nwaySelect_0n[10]);
  ND2 I937 (nwayMuxOut_10n[13], inp_10d[13], nwaySelect_0n[10]);
  ND2 I938 (nwayMuxOut_10n[14], inp_10d[14], nwaySelect_0n[10]);
  ND2 I939 (nwayMuxOut_10n[15], inp_10d[15], nwaySelect_0n[10]);
  ND2 I940 (nwayMuxOut_10n[16], inp_10d[16], nwaySelect_0n[10]);
  ND2 I941 (nwayMuxOut_10n[17], inp_10d[17], nwaySelect_0n[10]);
  ND2 I942 (nwayMuxOut_10n[18], inp_10d[18], nwaySelect_0n[10]);
  ND2 I943 (nwayMuxOut_10n[19], inp_10d[19], nwaySelect_0n[10]);
  ND2 I944 (nwayMuxOut_10n[20], inp_10d[20], nwaySelect_0n[10]);
  ND2 I945 (nwayMuxOut_10n[21], inp_10d[21], nwaySelect_0n[10]);
  ND2 I946 (nwayMuxOut_10n[22], inp_10d[22], nwaySelect_0n[10]);
  ND2 I947 (nwayMuxOut_10n[23], inp_10d[23], nwaySelect_0n[10]);
  ND2 I948 (nwayMuxOut_10n[24], inp_10d[24], nwaySelect_0n[10]);
  ND2 I949 (nwayMuxOut_10n[25], inp_10d[25], nwaySelect_0n[10]);
  ND2 I950 (nwayMuxOut_10n[26], inp_10d[26], nwaySelect_0n[10]);
  ND2 I951 (nwayMuxOut_10n[27], inp_10d[27], nwaySelect_0n[10]);
  ND2 I952 (nwayMuxOut_10n[28], inp_10d[28], nwaySelect_0n[10]);
  ND2 I953 (nwayMuxOut_10n[29], inp_10d[29], nwaySelect_0n[10]);
  ND2 I954 (nwayMuxOut_10n[30], inp_10d[30], nwaySelect_0n[10]);
  ND2 I955 (nwayMuxOut_10n[31], inp_10d[31], nwaySelect_0n[10]);
  ND2 I956 (nwayMuxOut_10n[32], inp_10d[32], nwaySelect_0n[10]);
  ND2 I957 (nwayMuxOut_11n[0], inp_11d[0], nwaySelect_0n[11]);
  ND2 I958 (nwayMuxOut_11n[1], inp_11d[1], nwaySelect_0n[11]);
  ND2 I959 (nwayMuxOut_11n[2], inp_11d[2], nwaySelect_0n[11]);
  ND2 I960 (nwayMuxOut_11n[3], inp_11d[3], nwaySelect_0n[11]);
  ND2 I961 (nwayMuxOut_11n[4], inp_11d[4], nwaySelect_0n[11]);
  ND2 I962 (nwayMuxOut_11n[5], inp_11d[5], nwaySelect_0n[11]);
  ND2 I963 (nwayMuxOut_11n[6], inp_11d[6], nwaySelect_0n[11]);
  ND2 I964 (nwayMuxOut_11n[7], inp_11d[7], nwaySelect_0n[11]);
  ND2 I965 (nwayMuxOut_11n[8], inp_11d[8], nwaySelect_0n[11]);
  ND2 I966 (nwayMuxOut_11n[9], inp_11d[9], nwaySelect_0n[11]);
  ND2 I967 (nwayMuxOut_11n[10], inp_11d[10], nwaySelect_0n[11]);
  ND2 I968 (nwayMuxOut_11n[11], inp_11d[11], nwaySelect_0n[11]);
  ND2 I969 (nwayMuxOut_11n[12], inp_11d[12], nwaySelect_0n[11]);
  ND2 I970 (nwayMuxOut_11n[13], inp_11d[13], nwaySelect_0n[11]);
  ND2 I971 (nwayMuxOut_11n[14], inp_11d[14], nwaySelect_0n[11]);
  ND2 I972 (nwayMuxOut_11n[15], inp_11d[15], nwaySelect_0n[11]);
  ND2 I973 (nwayMuxOut_11n[16], inp_11d[16], nwaySelect_0n[11]);
  ND2 I974 (nwayMuxOut_11n[17], inp_11d[17], nwaySelect_0n[11]);
  ND2 I975 (nwayMuxOut_11n[18], inp_11d[18], nwaySelect_0n[11]);
  ND2 I976 (nwayMuxOut_11n[19], inp_11d[19], nwaySelect_0n[11]);
  ND2 I977 (nwayMuxOut_11n[20], inp_11d[20], nwaySelect_0n[11]);
  ND2 I978 (nwayMuxOut_11n[21], inp_11d[21], nwaySelect_0n[11]);
  ND2 I979 (nwayMuxOut_11n[22], inp_11d[22], nwaySelect_0n[11]);
  ND2 I980 (nwayMuxOut_11n[23], inp_11d[23], nwaySelect_0n[11]);
  ND2 I981 (nwayMuxOut_11n[24], inp_11d[24], nwaySelect_0n[11]);
  ND2 I982 (nwayMuxOut_11n[25], inp_11d[25], nwaySelect_0n[11]);
  ND2 I983 (nwayMuxOut_11n[26], inp_11d[26], nwaySelect_0n[11]);
  ND2 I984 (nwayMuxOut_11n[27], inp_11d[27], nwaySelect_0n[11]);
  ND2 I985 (nwayMuxOut_11n[28], inp_11d[28], nwaySelect_0n[11]);
  ND2 I986 (nwayMuxOut_11n[29], inp_11d[29], nwaySelect_0n[11]);
  ND2 I987 (nwayMuxOut_11n[30], inp_11d[30], nwaySelect_0n[11]);
  ND2 I988 (nwayMuxOut_11n[31], inp_11d[31], nwaySelect_0n[11]);
  ND2 I989 (nwayMuxOut_11n[32], inp_11d[32], nwaySelect_0n[11]);
  ND2 I990 (nwayMuxOut_12n[0], inp_12d[0], nwaySelect_0n[12]);
  ND2 I991 (nwayMuxOut_12n[1], inp_12d[1], nwaySelect_0n[12]);
  ND2 I992 (nwayMuxOut_12n[2], inp_12d[2], nwaySelect_0n[12]);
  ND2 I993 (nwayMuxOut_12n[3], inp_12d[3], nwaySelect_0n[12]);
  ND2 I994 (nwayMuxOut_12n[4], inp_12d[4], nwaySelect_0n[12]);
  ND2 I995 (nwayMuxOut_12n[5], inp_12d[5], nwaySelect_0n[12]);
  ND2 I996 (nwayMuxOut_12n[6], inp_12d[6], nwaySelect_0n[12]);
  ND2 I997 (nwayMuxOut_12n[7], inp_12d[7], nwaySelect_0n[12]);
  ND2 I998 (nwayMuxOut_12n[8], inp_12d[8], nwaySelect_0n[12]);
  ND2 I999 (nwayMuxOut_12n[9], inp_12d[9], nwaySelect_0n[12]);
  ND2 I1000 (nwayMuxOut_12n[10], inp_12d[10], nwaySelect_0n[12]);
  ND2 I1001 (nwayMuxOut_12n[11], inp_12d[11], nwaySelect_0n[12]);
  ND2 I1002 (nwayMuxOut_12n[12], inp_12d[12], nwaySelect_0n[12]);
  ND2 I1003 (nwayMuxOut_12n[13], inp_12d[13], nwaySelect_0n[12]);
  ND2 I1004 (nwayMuxOut_12n[14], inp_12d[14], nwaySelect_0n[12]);
  ND2 I1005 (nwayMuxOut_12n[15], inp_12d[15], nwaySelect_0n[12]);
  ND2 I1006 (nwayMuxOut_12n[16], inp_12d[16], nwaySelect_0n[12]);
  ND2 I1007 (nwayMuxOut_12n[17], inp_12d[17], nwaySelect_0n[12]);
  ND2 I1008 (nwayMuxOut_12n[18], inp_12d[18], nwaySelect_0n[12]);
  ND2 I1009 (nwayMuxOut_12n[19], inp_12d[19], nwaySelect_0n[12]);
  ND2 I1010 (nwayMuxOut_12n[20], inp_12d[20], nwaySelect_0n[12]);
  ND2 I1011 (nwayMuxOut_12n[21], inp_12d[21], nwaySelect_0n[12]);
  ND2 I1012 (nwayMuxOut_12n[22], inp_12d[22], nwaySelect_0n[12]);
  ND2 I1013 (nwayMuxOut_12n[23], inp_12d[23], nwaySelect_0n[12]);
  ND2 I1014 (nwayMuxOut_12n[24], inp_12d[24], nwaySelect_0n[12]);
  ND2 I1015 (nwayMuxOut_12n[25], inp_12d[25], nwaySelect_0n[12]);
  ND2 I1016 (nwayMuxOut_12n[26], inp_12d[26], nwaySelect_0n[12]);
  ND2 I1017 (nwayMuxOut_12n[27], inp_12d[27], nwaySelect_0n[12]);
  ND2 I1018 (nwayMuxOut_12n[28], inp_12d[28], nwaySelect_0n[12]);
  ND2 I1019 (nwayMuxOut_12n[29], inp_12d[29], nwaySelect_0n[12]);
  ND2 I1020 (nwayMuxOut_12n[30], inp_12d[30], nwaySelect_0n[12]);
  ND2 I1021 (nwayMuxOut_12n[31], inp_12d[31], nwaySelect_0n[12]);
  ND2 I1022 (nwayMuxOut_12n[32], inp_12d[32], nwaySelect_0n[12]);
  ND2 I1023 (nwayMuxOut_13n[0], inp_13d[0], nwaySelect_0n[13]);
  ND2 I1024 (nwayMuxOut_13n[1], inp_13d[1], nwaySelect_0n[13]);
  ND2 I1025 (nwayMuxOut_13n[2], inp_13d[2], nwaySelect_0n[13]);
  ND2 I1026 (nwayMuxOut_13n[3], inp_13d[3], nwaySelect_0n[13]);
  ND2 I1027 (nwayMuxOut_13n[4], inp_13d[4], nwaySelect_0n[13]);
  ND2 I1028 (nwayMuxOut_13n[5], inp_13d[5], nwaySelect_0n[13]);
  ND2 I1029 (nwayMuxOut_13n[6], inp_13d[6], nwaySelect_0n[13]);
  ND2 I1030 (nwayMuxOut_13n[7], inp_13d[7], nwaySelect_0n[13]);
  ND2 I1031 (nwayMuxOut_13n[8], inp_13d[8], nwaySelect_0n[13]);
  ND2 I1032 (nwayMuxOut_13n[9], inp_13d[9], nwaySelect_0n[13]);
  ND2 I1033 (nwayMuxOut_13n[10], inp_13d[10], nwaySelect_0n[13]);
  ND2 I1034 (nwayMuxOut_13n[11], inp_13d[11], nwaySelect_0n[13]);
  ND2 I1035 (nwayMuxOut_13n[12], inp_13d[12], nwaySelect_0n[13]);
  ND2 I1036 (nwayMuxOut_13n[13], inp_13d[13], nwaySelect_0n[13]);
  ND2 I1037 (nwayMuxOut_13n[14], inp_13d[14], nwaySelect_0n[13]);
  ND2 I1038 (nwayMuxOut_13n[15], inp_13d[15], nwaySelect_0n[13]);
  ND2 I1039 (nwayMuxOut_13n[16], inp_13d[16], nwaySelect_0n[13]);
  ND2 I1040 (nwayMuxOut_13n[17], inp_13d[17], nwaySelect_0n[13]);
  ND2 I1041 (nwayMuxOut_13n[18], inp_13d[18], nwaySelect_0n[13]);
  ND2 I1042 (nwayMuxOut_13n[19], inp_13d[19], nwaySelect_0n[13]);
  ND2 I1043 (nwayMuxOut_13n[20], inp_13d[20], nwaySelect_0n[13]);
  ND2 I1044 (nwayMuxOut_13n[21], inp_13d[21], nwaySelect_0n[13]);
  ND2 I1045 (nwayMuxOut_13n[22], inp_13d[22], nwaySelect_0n[13]);
  ND2 I1046 (nwayMuxOut_13n[23], inp_13d[23], nwaySelect_0n[13]);
  ND2 I1047 (nwayMuxOut_13n[24], inp_13d[24], nwaySelect_0n[13]);
  ND2 I1048 (nwayMuxOut_13n[25], inp_13d[25], nwaySelect_0n[13]);
  ND2 I1049 (nwayMuxOut_13n[26], inp_13d[26], nwaySelect_0n[13]);
  ND2 I1050 (nwayMuxOut_13n[27], inp_13d[27], nwaySelect_0n[13]);
  ND2 I1051 (nwayMuxOut_13n[28], inp_13d[28], nwaySelect_0n[13]);
  ND2 I1052 (nwayMuxOut_13n[29], inp_13d[29], nwaySelect_0n[13]);
  ND2 I1053 (nwayMuxOut_13n[30], inp_13d[30], nwaySelect_0n[13]);
  ND2 I1054 (nwayMuxOut_13n[31], inp_13d[31], nwaySelect_0n[13]);
  ND2 I1055 (nwayMuxOut_13n[32], inp_13d[32], nwaySelect_0n[13]);
  ND2 I1056 (nwayMuxOut_14n[0], inp_14d[0], nwaySelect_0n[14]);
  ND2 I1057 (nwayMuxOut_14n[1], inp_14d[1], nwaySelect_0n[14]);
  ND2 I1058 (nwayMuxOut_14n[2], inp_14d[2], nwaySelect_0n[14]);
  ND2 I1059 (nwayMuxOut_14n[3], inp_14d[3], nwaySelect_0n[14]);
  ND2 I1060 (nwayMuxOut_14n[4], inp_14d[4], nwaySelect_0n[14]);
  ND2 I1061 (nwayMuxOut_14n[5], inp_14d[5], nwaySelect_0n[14]);
  ND2 I1062 (nwayMuxOut_14n[6], inp_14d[6], nwaySelect_0n[14]);
  ND2 I1063 (nwayMuxOut_14n[7], inp_14d[7], nwaySelect_0n[14]);
  ND2 I1064 (nwayMuxOut_14n[8], inp_14d[8], nwaySelect_0n[14]);
  ND2 I1065 (nwayMuxOut_14n[9], inp_14d[9], nwaySelect_0n[14]);
  ND2 I1066 (nwayMuxOut_14n[10], inp_14d[10], nwaySelect_0n[14]);
  ND2 I1067 (nwayMuxOut_14n[11], inp_14d[11], nwaySelect_0n[14]);
  ND2 I1068 (nwayMuxOut_14n[12], inp_14d[12], nwaySelect_0n[14]);
  ND2 I1069 (nwayMuxOut_14n[13], inp_14d[13], nwaySelect_0n[14]);
  ND2 I1070 (nwayMuxOut_14n[14], inp_14d[14], nwaySelect_0n[14]);
  ND2 I1071 (nwayMuxOut_14n[15], inp_14d[15], nwaySelect_0n[14]);
  ND2 I1072 (nwayMuxOut_14n[16], inp_14d[16], nwaySelect_0n[14]);
  ND2 I1073 (nwayMuxOut_14n[17], inp_14d[17], nwaySelect_0n[14]);
  ND2 I1074 (nwayMuxOut_14n[18], inp_14d[18], nwaySelect_0n[14]);
  ND2 I1075 (nwayMuxOut_14n[19], inp_14d[19], nwaySelect_0n[14]);
  ND2 I1076 (nwayMuxOut_14n[20], inp_14d[20], nwaySelect_0n[14]);
  ND2 I1077 (nwayMuxOut_14n[21], inp_14d[21], nwaySelect_0n[14]);
  ND2 I1078 (nwayMuxOut_14n[22], inp_14d[22], nwaySelect_0n[14]);
  ND2 I1079 (nwayMuxOut_14n[23], inp_14d[23], nwaySelect_0n[14]);
  ND2 I1080 (nwayMuxOut_14n[24], inp_14d[24], nwaySelect_0n[14]);
  ND2 I1081 (nwayMuxOut_14n[25], inp_14d[25], nwaySelect_0n[14]);
  ND2 I1082 (nwayMuxOut_14n[26], inp_14d[26], nwaySelect_0n[14]);
  ND2 I1083 (nwayMuxOut_14n[27], inp_14d[27], nwaySelect_0n[14]);
  ND2 I1084 (nwayMuxOut_14n[28], inp_14d[28], nwaySelect_0n[14]);
  ND2 I1085 (nwayMuxOut_14n[29], inp_14d[29], nwaySelect_0n[14]);
  ND2 I1086 (nwayMuxOut_14n[30], inp_14d[30], nwaySelect_0n[14]);
  ND2 I1087 (nwayMuxOut_14n[31], inp_14d[31], nwaySelect_0n[14]);
  ND2 I1088 (nwayMuxOut_14n[32], inp_14d[32], nwaySelect_0n[14]);
  ND2 I1089 (nwayMuxOut_15n[0], inp_15d[0], nwaySelect_0n[15]);
  ND2 I1090 (nwayMuxOut_15n[1], inp_15d[1], nwaySelect_0n[15]);
  ND2 I1091 (nwayMuxOut_15n[2], inp_15d[2], nwaySelect_0n[15]);
  ND2 I1092 (nwayMuxOut_15n[3], inp_15d[3], nwaySelect_0n[15]);
  ND2 I1093 (nwayMuxOut_15n[4], inp_15d[4], nwaySelect_0n[15]);
  ND2 I1094 (nwayMuxOut_15n[5], inp_15d[5], nwaySelect_0n[15]);
  ND2 I1095 (nwayMuxOut_15n[6], inp_15d[6], nwaySelect_0n[15]);
  ND2 I1096 (nwayMuxOut_15n[7], inp_15d[7], nwaySelect_0n[15]);
  ND2 I1097 (nwayMuxOut_15n[8], inp_15d[8], nwaySelect_0n[15]);
  ND2 I1098 (nwayMuxOut_15n[9], inp_15d[9], nwaySelect_0n[15]);
  ND2 I1099 (nwayMuxOut_15n[10], inp_15d[10], nwaySelect_0n[15]);
  ND2 I1100 (nwayMuxOut_15n[11], inp_15d[11], nwaySelect_0n[15]);
  ND2 I1101 (nwayMuxOut_15n[12], inp_15d[12], nwaySelect_0n[15]);
  ND2 I1102 (nwayMuxOut_15n[13], inp_15d[13], nwaySelect_0n[15]);
  ND2 I1103 (nwayMuxOut_15n[14], inp_15d[14], nwaySelect_0n[15]);
  ND2 I1104 (nwayMuxOut_15n[15], inp_15d[15], nwaySelect_0n[15]);
  ND2 I1105 (nwayMuxOut_15n[16], inp_15d[16], nwaySelect_0n[15]);
  ND2 I1106 (nwayMuxOut_15n[17], inp_15d[17], nwaySelect_0n[15]);
  ND2 I1107 (nwayMuxOut_15n[18], inp_15d[18], nwaySelect_0n[15]);
  ND2 I1108 (nwayMuxOut_15n[19], inp_15d[19], nwaySelect_0n[15]);
  ND2 I1109 (nwayMuxOut_15n[20], inp_15d[20], nwaySelect_0n[15]);
  ND2 I1110 (nwayMuxOut_15n[21], inp_15d[21], nwaySelect_0n[15]);
  ND2 I1111 (nwayMuxOut_15n[22], inp_15d[22], nwaySelect_0n[15]);
  ND2 I1112 (nwayMuxOut_15n[23], inp_15d[23], nwaySelect_0n[15]);
  ND2 I1113 (nwayMuxOut_15n[24], inp_15d[24], nwaySelect_0n[15]);
  ND2 I1114 (nwayMuxOut_15n[25], inp_15d[25], nwaySelect_0n[15]);
  ND2 I1115 (nwayMuxOut_15n[26], inp_15d[26], nwaySelect_0n[15]);
  ND2 I1116 (nwayMuxOut_15n[27], inp_15d[27], nwaySelect_0n[15]);
  ND2 I1117 (nwayMuxOut_15n[28], inp_15d[28], nwaySelect_0n[15]);
  ND2 I1118 (nwayMuxOut_15n[29], inp_15d[29], nwaySelect_0n[15]);
  ND2 I1119 (nwayMuxOut_15n[30], inp_15d[30], nwaySelect_0n[15]);
  ND2 I1120 (nwayMuxOut_15n[31], inp_15d[31], nwaySelect_0n[15]);
  ND2 I1121 (nwayMuxOut_15n[32], inp_15d[32], nwaySelect_0n[15]);
  ND2 I1122 (nwayMuxOut_16n[0], inp_16d[0], nwaySelect_0n[16]);
  ND2 I1123 (nwayMuxOut_16n[1], inp_16d[1], nwaySelect_0n[16]);
  ND2 I1124 (nwayMuxOut_16n[2], inp_16d[2], nwaySelect_0n[16]);
  ND2 I1125 (nwayMuxOut_16n[3], inp_16d[3], nwaySelect_0n[16]);
  ND2 I1126 (nwayMuxOut_16n[4], inp_16d[4], nwaySelect_0n[16]);
  ND2 I1127 (nwayMuxOut_16n[5], inp_16d[5], nwaySelect_0n[16]);
  ND2 I1128 (nwayMuxOut_16n[6], inp_16d[6], nwaySelect_0n[16]);
  ND2 I1129 (nwayMuxOut_16n[7], inp_16d[7], nwaySelect_0n[16]);
  ND2 I1130 (nwayMuxOut_16n[8], inp_16d[8], nwaySelect_0n[16]);
  ND2 I1131 (nwayMuxOut_16n[9], inp_16d[9], nwaySelect_0n[16]);
  ND2 I1132 (nwayMuxOut_16n[10], inp_16d[10], nwaySelect_0n[16]);
  ND2 I1133 (nwayMuxOut_16n[11], inp_16d[11], nwaySelect_0n[16]);
  ND2 I1134 (nwayMuxOut_16n[12], inp_16d[12], nwaySelect_0n[16]);
  ND2 I1135 (nwayMuxOut_16n[13], inp_16d[13], nwaySelect_0n[16]);
  ND2 I1136 (nwayMuxOut_16n[14], inp_16d[14], nwaySelect_0n[16]);
  ND2 I1137 (nwayMuxOut_16n[15], inp_16d[15], nwaySelect_0n[16]);
  ND2 I1138 (nwayMuxOut_16n[16], inp_16d[16], nwaySelect_0n[16]);
  ND2 I1139 (nwayMuxOut_16n[17], inp_16d[17], nwaySelect_0n[16]);
  ND2 I1140 (nwayMuxOut_16n[18], inp_16d[18], nwaySelect_0n[16]);
  ND2 I1141 (nwayMuxOut_16n[19], inp_16d[19], nwaySelect_0n[16]);
  ND2 I1142 (nwayMuxOut_16n[20], inp_16d[20], nwaySelect_0n[16]);
  ND2 I1143 (nwayMuxOut_16n[21], inp_16d[21], nwaySelect_0n[16]);
  ND2 I1144 (nwayMuxOut_16n[22], inp_16d[22], nwaySelect_0n[16]);
  ND2 I1145 (nwayMuxOut_16n[23], inp_16d[23], nwaySelect_0n[16]);
  ND2 I1146 (nwayMuxOut_16n[24], inp_16d[24], nwaySelect_0n[16]);
  ND2 I1147 (nwayMuxOut_16n[25], inp_16d[25], nwaySelect_0n[16]);
  ND2 I1148 (nwayMuxOut_16n[26], inp_16d[26], nwaySelect_0n[16]);
  ND2 I1149 (nwayMuxOut_16n[27], inp_16d[27], nwaySelect_0n[16]);
  ND2 I1150 (nwayMuxOut_16n[28], inp_16d[28], nwaySelect_0n[16]);
  ND2 I1151 (nwayMuxOut_16n[29], inp_16d[29], nwaySelect_0n[16]);
  ND2 I1152 (nwayMuxOut_16n[30], inp_16d[30], nwaySelect_0n[16]);
  ND2 I1153 (nwayMuxOut_16n[31], inp_16d[31], nwaySelect_0n[16]);
  ND2 I1154 (nwayMuxOut_16n[32], inp_16d[32], nwaySelect_0n[16]);
  ND2 I1155 (nwayMuxOut_17n[0], inp_17d[0], nwaySelect_0n[17]);
  ND2 I1156 (nwayMuxOut_17n[1], inp_17d[1], nwaySelect_0n[17]);
  ND2 I1157 (nwayMuxOut_17n[2], inp_17d[2], nwaySelect_0n[17]);
  ND2 I1158 (nwayMuxOut_17n[3], inp_17d[3], nwaySelect_0n[17]);
  ND2 I1159 (nwayMuxOut_17n[4], inp_17d[4], nwaySelect_0n[17]);
  ND2 I1160 (nwayMuxOut_17n[5], inp_17d[5], nwaySelect_0n[17]);
  ND2 I1161 (nwayMuxOut_17n[6], inp_17d[6], nwaySelect_0n[17]);
  ND2 I1162 (nwayMuxOut_17n[7], inp_17d[7], nwaySelect_0n[17]);
  ND2 I1163 (nwayMuxOut_17n[8], inp_17d[8], nwaySelect_0n[17]);
  ND2 I1164 (nwayMuxOut_17n[9], inp_17d[9], nwaySelect_0n[17]);
  ND2 I1165 (nwayMuxOut_17n[10], inp_17d[10], nwaySelect_0n[17]);
  ND2 I1166 (nwayMuxOut_17n[11], inp_17d[11], nwaySelect_0n[17]);
  ND2 I1167 (nwayMuxOut_17n[12], inp_17d[12], nwaySelect_0n[17]);
  ND2 I1168 (nwayMuxOut_17n[13], inp_17d[13], nwaySelect_0n[17]);
  ND2 I1169 (nwayMuxOut_17n[14], inp_17d[14], nwaySelect_0n[17]);
  ND2 I1170 (nwayMuxOut_17n[15], inp_17d[15], nwaySelect_0n[17]);
  ND2 I1171 (nwayMuxOut_17n[16], inp_17d[16], nwaySelect_0n[17]);
  ND2 I1172 (nwayMuxOut_17n[17], inp_17d[17], nwaySelect_0n[17]);
  ND2 I1173 (nwayMuxOut_17n[18], inp_17d[18], nwaySelect_0n[17]);
  ND2 I1174 (nwayMuxOut_17n[19], inp_17d[19], nwaySelect_0n[17]);
  ND2 I1175 (nwayMuxOut_17n[20], inp_17d[20], nwaySelect_0n[17]);
  ND2 I1176 (nwayMuxOut_17n[21], inp_17d[21], nwaySelect_0n[17]);
  ND2 I1177 (nwayMuxOut_17n[22], inp_17d[22], nwaySelect_0n[17]);
  ND2 I1178 (nwayMuxOut_17n[23], inp_17d[23], nwaySelect_0n[17]);
  ND2 I1179 (nwayMuxOut_17n[24], inp_17d[24], nwaySelect_0n[17]);
  ND2 I1180 (nwayMuxOut_17n[25], inp_17d[25], nwaySelect_0n[17]);
  ND2 I1181 (nwayMuxOut_17n[26], inp_17d[26], nwaySelect_0n[17]);
  ND2 I1182 (nwayMuxOut_17n[27], inp_17d[27], nwaySelect_0n[17]);
  ND2 I1183 (nwayMuxOut_17n[28], inp_17d[28], nwaySelect_0n[17]);
  ND2 I1184 (nwayMuxOut_17n[29], inp_17d[29], nwaySelect_0n[17]);
  ND2 I1185 (nwayMuxOut_17n[30], inp_17d[30], nwaySelect_0n[17]);
  ND2 I1186 (nwayMuxOut_17n[31], inp_17d[31], nwaySelect_0n[17]);
  ND2 I1187 (nwayMuxOut_17n[32], inp_17d[32], nwaySelect_0n[17]);
  ND2 I1188 (nwayMuxOut_18n[0], inp_18d[0], nwaySelect_0n[18]);
  ND2 I1189 (nwayMuxOut_18n[1], inp_18d[1], nwaySelect_0n[18]);
  ND2 I1190 (nwayMuxOut_18n[2], inp_18d[2], nwaySelect_0n[18]);
  ND2 I1191 (nwayMuxOut_18n[3], inp_18d[3], nwaySelect_0n[18]);
  ND2 I1192 (nwayMuxOut_18n[4], inp_18d[4], nwaySelect_0n[18]);
  ND2 I1193 (nwayMuxOut_18n[5], inp_18d[5], nwaySelect_0n[18]);
  ND2 I1194 (nwayMuxOut_18n[6], inp_18d[6], nwaySelect_0n[18]);
  ND2 I1195 (nwayMuxOut_18n[7], inp_18d[7], nwaySelect_0n[18]);
  ND2 I1196 (nwayMuxOut_18n[8], inp_18d[8], nwaySelect_0n[18]);
  ND2 I1197 (nwayMuxOut_18n[9], inp_18d[9], nwaySelect_0n[18]);
  ND2 I1198 (nwayMuxOut_18n[10], inp_18d[10], nwaySelect_0n[18]);
  ND2 I1199 (nwayMuxOut_18n[11], inp_18d[11], nwaySelect_0n[18]);
  ND2 I1200 (nwayMuxOut_18n[12], inp_18d[12], nwaySelect_0n[18]);
  ND2 I1201 (nwayMuxOut_18n[13], inp_18d[13], nwaySelect_0n[18]);
  ND2 I1202 (nwayMuxOut_18n[14], inp_18d[14], nwaySelect_0n[18]);
  ND2 I1203 (nwayMuxOut_18n[15], inp_18d[15], nwaySelect_0n[18]);
  ND2 I1204 (nwayMuxOut_18n[16], inp_18d[16], nwaySelect_0n[18]);
  ND2 I1205 (nwayMuxOut_18n[17], inp_18d[17], nwaySelect_0n[18]);
  ND2 I1206 (nwayMuxOut_18n[18], inp_18d[18], nwaySelect_0n[18]);
  ND2 I1207 (nwayMuxOut_18n[19], inp_18d[19], nwaySelect_0n[18]);
  ND2 I1208 (nwayMuxOut_18n[20], inp_18d[20], nwaySelect_0n[18]);
  ND2 I1209 (nwayMuxOut_18n[21], inp_18d[21], nwaySelect_0n[18]);
  ND2 I1210 (nwayMuxOut_18n[22], inp_18d[22], nwaySelect_0n[18]);
  ND2 I1211 (nwayMuxOut_18n[23], inp_18d[23], nwaySelect_0n[18]);
  ND2 I1212 (nwayMuxOut_18n[24], inp_18d[24], nwaySelect_0n[18]);
  ND2 I1213 (nwayMuxOut_18n[25], inp_18d[25], nwaySelect_0n[18]);
  ND2 I1214 (nwayMuxOut_18n[26], inp_18d[26], nwaySelect_0n[18]);
  ND2 I1215 (nwayMuxOut_18n[27], inp_18d[27], nwaySelect_0n[18]);
  ND2 I1216 (nwayMuxOut_18n[28], inp_18d[28], nwaySelect_0n[18]);
  ND2 I1217 (nwayMuxOut_18n[29], inp_18d[29], nwaySelect_0n[18]);
  ND2 I1218 (nwayMuxOut_18n[30], inp_18d[30], nwaySelect_0n[18]);
  ND2 I1219 (nwayMuxOut_18n[31], inp_18d[31], nwaySelect_0n[18]);
  ND2 I1220 (nwayMuxOut_18n[32], inp_18d[32], nwaySelect_0n[18]);
  ND2 I1221 (nwayMuxOut_19n[0], inp_19d[0], nwaySelect_0n[19]);
  ND2 I1222 (nwayMuxOut_19n[1], inp_19d[1], nwaySelect_0n[19]);
  ND2 I1223 (nwayMuxOut_19n[2], inp_19d[2], nwaySelect_0n[19]);
  ND2 I1224 (nwayMuxOut_19n[3], inp_19d[3], nwaySelect_0n[19]);
  ND2 I1225 (nwayMuxOut_19n[4], inp_19d[4], nwaySelect_0n[19]);
  ND2 I1226 (nwayMuxOut_19n[5], inp_19d[5], nwaySelect_0n[19]);
  ND2 I1227 (nwayMuxOut_19n[6], inp_19d[6], nwaySelect_0n[19]);
  ND2 I1228 (nwayMuxOut_19n[7], inp_19d[7], nwaySelect_0n[19]);
  ND2 I1229 (nwayMuxOut_19n[8], inp_19d[8], nwaySelect_0n[19]);
  ND2 I1230 (nwayMuxOut_19n[9], inp_19d[9], nwaySelect_0n[19]);
  ND2 I1231 (nwayMuxOut_19n[10], inp_19d[10], nwaySelect_0n[19]);
  ND2 I1232 (nwayMuxOut_19n[11], inp_19d[11], nwaySelect_0n[19]);
  ND2 I1233 (nwayMuxOut_19n[12], inp_19d[12], nwaySelect_0n[19]);
  ND2 I1234 (nwayMuxOut_19n[13], inp_19d[13], nwaySelect_0n[19]);
  ND2 I1235 (nwayMuxOut_19n[14], inp_19d[14], nwaySelect_0n[19]);
  ND2 I1236 (nwayMuxOut_19n[15], inp_19d[15], nwaySelect_0n[19]);
  ND2 I1237 (nwayMuxOut_19n[16], inp_19d[16], nwaySelect_0n[19]);
  ND2 I1238 (nwayMuxOut_19n[17], inp_19d[17], nwaySelect_0n[19]);
  ND2 I1239 (nwayMuxOut_19n[18], inp_19d[18], nwaySelect_0n[19]);
  ND2 I1240 (nwayMuxOut_19n[19], inp_19d[19], nwaySelect_0n[19]);
  ND2 I1241 (nwayMuxOut_19n[20], inp_19d[20], nwaySelect_0n[19]);
  ND2 I1242 (nwayMuxOut_19n[21], inp_19d[21], nwaySelect_0n[19]);
  ND2 I1243 (nwayMuxOut_19n[22], inp_19d[22], nwaySelect_0n[19]);
  ND2 I1244 (nwayMuxOut_19n[23], inp_19d[23], nwaySelect_0n[19]);
  ND2 I1245 (nwayMuxOut_19n[24], inp_19d[24], nwaySelect_0n[19]);
  ND2 I1246 (nwayMuxOut_19n[25], inp_19d[25], nwaySelect_0n[19]);
  ND2 I1247 (nwayMuxOut_19n[26], inp_19d[26], nwaySelect_0n[19]);
  ND2 I1248 (nwayMuxOut_19n[27], inp_19d[27], nwaySelect_0n[19]);
  ND2 I1249 (nwayMuxOut_19n[28], inp_19d[28], nwaySelect_0n[19]);
  ND2 I1250 (nwayMuxOut_19n[29], inp_19d[29], nwaySelect_0n[19]);
  ND2 I1251 (nwayMuxOut_19n[30], inp_19d[30], nwaySelect_0n[19]);
  ND2 I1252 (nwayMuxOut_19n[31], inp_19d[31], nwaySelect_0n[19]);
  ND2 I1253 (nwayMuxOut_19n[32], inp_19d[32], nwaySelect_0n[19]);
  ND2 I1254 (nwayMuxOut_20n[0], inp_20d[0], nwaySelect_0n[20]);
  ND2 I1255 (nwayMuxOut_20n[1], inp_20d[1], nwaySelect_0n[20]);
  ND2 I1256 (nwayMuxOut_20n[2], inp_20d[2], nwaySelect_0n[20]);
  ND2 I1257 (nwayMuxOut_20n[3], inp_20d[3], nwaySelect_0n[20]);
  ND2 I1258 (nwayMuxOut_20n[4], inp_20d[4], nwaySelect_0n[20]);
  ND2 I1259 (nwayMuxOut_20n[5], inp_20d[5], nwaySelect_0n[20]);
  ND2 I1260 (nwayMuxOut_20n[6], inp_20d[6], nwaySelect_0n[20]);
  ND2 I1261 (nwayMuxOut_20n[7], inp_20d[7], nwaySelect_0n[20]);
  ND2 I1262 (nwayMuxOut_20n[8], inp_20d[8], nwaySelect_0n[20]);
  ND2 I1263 (nwayMuxOut_20n[9], inp_20d[9], nwaySelect_0n[20]);
  ND2 I1264 (nwayMuxOut_20n[10], inp_20d[10], nwaySelect_0n[20]);
  ND2 I1265 (nwayMuxOut_20n[11], inp_20d[11], nwaySelect_0n[20]);
  ND2 I1266 (nwayMuxOut_20n[12], inp_20d[12], nwaySelect_0n[20]);
  ND2 I1267 (nwayMuxOut_20n[13], inp_20d[13], nwaySelect_0n[20]);
  ND2 I1268 (nwayMuxOut_20n[14], inp_20d[14], nwaySelect_0n[20]);
  ND2 I1269 (nwayMuxOut_20n[15], inp_20d[15], nwaySelect_0n[20]);
  ND2 I1270 (nwayMuxOut_20n[16], inp_20d[16], nwaySelect_0n[20]);
  ND2 I1271 (nwayMuxOut_20n[17], inp_20d[17], nwaySelect_0n[20]);
  ND2 I1272 (nwayMuxOut_20n[18], inp_20d[18], nwaySelect_0n[20]);
  ND2 I1273 (nwayMuxOut_20n[19], inp_20d[19], nwaySelect_0n[20]);
  ND2 I1274 (nwayMuxOut_20n[20], inp_20d[20], nwaySelect_0n[20]);
  ND2 I1275 (nwayMuxOut_20n[21], inp_20d[21], nwaySelect_0n[20]);
  ND2 I1276 (nwayMuxOut_20n[22], inp_20d[22], nwaySelect_0n[20]);
  ND2 I1277 (nwayMuxOut_20n[23], inp_20d[23], nwaySelect_0n[20]);
  ND2 I1278 (nwayMuxOut_20n[24], inp_20d[24], nwaySelect_0n[20]);
  ND2 I1279 (nwayMuxOut_20n[25], inp_20d[25], nwaySelect_0n[20]);
  ND2 I1280 (nwayMuxOut_20n[26], inp_20d[26], nwaySelect_0n[20]);
  ND2 I1281 (nwayMuxOut_20n[27], inp_20d[27], nwaySelect_0n[20]);
  ND2 I1282 (nwayMuxOut_20n[28], inp_20d[28], nwaySelect_0n[20]);
  ND2 I1283 (nwayMuxOut_20n[29], inp_20d[29], nwaySelect_0n[20]);
  ND2 I1284 (nwayMuxOut_20n[30], inp_20d[30], nwaySelect_0n[20]);
  ND2 I1285 (nwayMuxOut_20n[31], inp_20d[31], nwaySelect_0n[20]);
  ND2 I1286 (nwayMuxOut_20n[32], inp_20d[32], nwaySelect_0n[20]);
  ND2 I1287 (nwayMuxOut_21n[0], inp_21d[0], nwaySelect_0n[21]);
  ND2 I1288 (nwayMuxOut_21n[1], inp_21d[1], nwaySelect_0n[21]);
  ND2 I1289 (nwayMuxOut_21n[2], inp_21d[2], nwaySelect_0n[21]);
  ND2 I1290 (nwayMuxOut_21n[3], inp_21d[3], nwaySelect_0n[21]);
  ND2 I1291 (nwayMuxOut_21n[4], inp_21d[4], nwaySelect_0n[21]);
  ND2 I1292 (nwayMuxOut_21n[5], inp_21d[5], nwaySelect_0n[21]);
  ND2 I1293 (nwayMuxOut_21n[6], inp_21d[6], nwaySelect_0n[21]);
  ND2 I1294 (nwayMuxOut_21n[7], inp_21d[7], nwaySelect_0n[21]);
  ND2 I1295 (nwayMuxOut_21n[8], inp_21d[8], nwaySelect_0n[21]);
  ND2 I1296 (nwayMuxOut_21n[9], inp_21d[9], nwaySelect_0n[21]);
  ND2 I1297 (nwayMuxOut_21n[10], inp_21d[10], nwaySelect_0n[21]);
  ND2 I1298 (nwayMuxOut_21n[11], inp_21d[11], nwaySelect_0n[21]);
  ND2 I1299 (nwayMuxOut_21n[12], inp_21d[12], nwaySelect_0n[21]);
  ND2 I1300 (nwayMuxOut_21n[13], inp_21d[13], nwaySelect_0n[21]);
  ND2 I1301 (nwayMuxOut_21n[14], inp_21d[14], nwaySelect_0n[21]);
  ND2 I1302 (nwayMuxOut_21n[15], inp_21d[15], nwaySelect_0n[21]);
  ND2 I1303 (nwayMuxOut_21n[16], inp_21d[16], nwaySelect_0n[21]);
  ND2 I1304 (nwayMuxOut_21n[17], inp_21d[17], nwaySelect_0n[21]);
  ND2 I1305 (nwayMuxOut_21n[18], inp_21d[18], nwaySelect_0n[21]);
  ND2 I1306 (nwayMuxOut_21n[19], inp_21d[19], nwaySelect_0n[21]);
  ND2 I1307 (nwayMuxOut_21n[20], inp_21d[20], nwaySelect_0n[21]);
  ND2 I1308 (nwayMuxOut_21n[21], inp_21d[21], nwaySelect_0n[21]);
  ND2 I1309 (nwayMuxOut_21n[22], inp_21d[22], nwaySelect_0n[21]);
  ND2 I1310 (nwayMuxOut_21n[23], inp_21d[23], nwaySelect_0n[21]);
  ND2 I1311 (nwayMuxOut_21n[24], inp_21d[24], nwaySelect_0n[21]);
  ND2 I1312 (nwayMuxOut_21n[25], inp_21d[25], nwaySelect_0n[21]);
  ND2 I1313 (nwayMuxOut_21n[26], inp_21d[26], nwaySelect_0n[21]);
  ND2 I1314 (nwayMuxOut_21n[27], inp_21d[27], nwaySelect_0n[21]);
  ND2 I1315 (nwayMuxOut_21n[28], inp_21d[28], nwaySelect_0n[21]);
  ND2 I1316 (nwayMuxOut_21n[29], inp_21d[29], nwaySelect_0n[21]);
  ND2 I1317 (nwayMuxOut_21n[30], inp_21d[30], nwaySelect_0n[21]);
  ND2 I1318 (nwayMuxOut_21n[31], inp_21d[31], nwaySelect_0n[21]);
  ND2 I1319 (nwayMuxOut_21n[32], inp_21d[32], nwaySelect_0n[21]);
  ND2 I1320 (nwayMuxOut_22n[0], inp_22d[0], nwaySelect_0n[22]);
  ND2 I1321 (nwayMuxOut_22n[1], inp_22d[1], nwaySelect_0n[22]);
  ND2 I1322 (nwayMuxOut_22n[2], inp_22d[2], nwaySelect_0n[22]);
  ND2 I1323 (nwayMuxOut_22n[3], inp_22d[3], nwaySelect_0n[22]);
  ND2 I1324 (nwayMuxOut_22n[4], inp_22d[4], nwaySelect_0n[22]);
  ND2 I1325 (nwayMuxOut_22n[5], inp_22d[5], nwaySelect_0n[22]);
  ND2 I1326 (nwayMuxOut_22n[6], inp_22d[6], nwaySelect_0n[22]);
  ND2 I1327 (nwayMuxOut_22n[7], inp_22d[7], nwaySelect_0n[22]);
  ND2 I1328 (nwayMuxOut_22n[8], inp_22d[8], nwaySelect_0n[22]);
  ND2 I1329 (nwayMuxOut_22n[9], inp_22d[9], nwaySelect_0n[22]);
  ND2 I1330 (nwayMuxOut_22n[10], inp_22d[10], nwaySelect_0n[22]);
  ND2 I1331 (nwayMuxOut_22n[11], inp_22d[11], nwaySelect_0n[22]);
  ND2 I1332 (nwayMuxOut_22n[12], inp_22d[12], nwaySelect_0n[22]);
  ND2 I1333 (nwayMuxOut_22n[13], inp_22d[13], nwaySelect_0n[22]);
  ND2 I1334 (nwayMuxOut_22n[14], inp_22d[14], nwaySelect_0n[22]);
  ND2 I1335 (nwayMuxOut_22n[15], inp_22d[15], nwaySelect_0n[22]);
  ND2 I1336 (nwayMuxOut_22n[16], inp_22d[16], nwaySelect_0n[22]);
  ND2 I1337 (nwayMuxOut_22n[17], inp_22d[17], nwaySelect_0n[22]);
  ND2 I1338 (nwayMuxOut_22n[18], inp_22d[18], nwaySelect_0n[22]);
  ND2 I1339 (nwayMuxOut_22n[19], inp_22d[19], nwaySelect_0n[22]);
  ND2 I1340 (nwayMuxOut_22n[20], inp_22d[20], nwaySelect_0n[22]);
  ND2 I1341 (nwayMuxOut_22n[21], inp_22d[21], nwaySelect_0n[22]);
  ND2 I1342 (nwayMuxOut_22n[22], inp_22d[22], nwaySelect_0n[22]);
  ND2 I1343 (nwayMuxOut_22n[23], inp_22d[23], nwaySelect_0n[22]);
  ND2 I1344 (nwayMuxOut_22n[24], inp_22d[24], nwaySelect_0n[22]);
  ND2 I1345 (nwayMuxOut_22n[25], inp_22d[25], nwaySelect_0n[22]);
  ND2 I1346 (nwayMuxOut_22n[26], inp_22d[26], nwaySelect_0n[22]);
  ND2 I1347 (nwayMuxOut_22n[27], inp_22d[27], nwaySelect_0n[22]);
  ND2 I1348 (nwayMuxOut_22n[28], inp_22d[28], nwaySelect_0n[22]);
  ND2 I1349 (nwayMuxOut_22n[29], inp_22d[29], nwaySelect_0n[22]);
  ND2 I1350 (nwayMuxOut_22n[30], inp_22d[30], nwaySelect_0n[22]);
  ND2 I1351 (nwayMuxOut_22n[31], inp_22d[31], nwaySelect_0n[22]);
  ND2 I1352 (nwayMuxOut_22n[32], inp_22d[32], nwaySelect_0n[22]);
  ND2 I1353 (nwayMuxOut_23n[0], inp_23d[0], nwaySelect_0n[23]);
  ND2 I1354 (nwayMuxOut_23n[1], inp_23d[1], nwaySelect_0n[23]);
  ND2 I1355 (nwayMuxOut_23n[2], inp_23d[2], nwaySelect_0n[23]);
  ND2 I1356 (nwayMuxOut_23n[3], inp_23d[3], nwaySelect_0n[23]);
  ND2 I1357 (nwayMuxOut_23n[4], inp_23d[4], nwaySelect_0n[23]);
  ND2 I1358 (nwayMuxOut_23n[5], inp_23d[5], nwaySelect_0n[23]);
  ND2 I1359 (nwayMuxOut_23n[6], inp_23d[6], nwaySelect_0n[23]);
  ND2 I1360 (nwayMuxOut_23n[7], inp_23d[7], nwaySelect_0n[23]);
  ND2 I1361 (nwayMuxOut_23n[8], inp_23d[8], nwaySelect_0n[23]);
  ND2 I1362 (nwayMuxOut_23n[9], inp_23d[9], nwaySelect_0n[23]);
  ND2 I1363 (nwayMuxOut_23n[10], inp_23d[10], nwaySelect_0n[23]);
  ND2 I1364 (nwayMuxOut_23n[11], inp_23d[11], nwaySelect_0n[23]);
  ND2 I1365 (nwayMuxOut_23n[12], inp_23d[12], nwaySelect_0n[23]);
  ND2 I1366 (nwayMuxOut_23n[13], inp_23d[13], nwaySelect_0n[23]);
  ND2 I1367 (nwayMuxOut_23n[14], inp_23d[14], nwaySelect_0n[23]);
  ND2 I1368 (nwayMuxOut_23n[15], inp_23d[15], nwaySelect_0n[23]);
  ND2 I1369 (nwayMuxOut_23n[16], inp_23d[16], nwaySelect_0n[23]);
  ND2 I1370 (nwayMuxOut_23n[17], inp_23d[17], nwaySelect_0n[23]);
  ND2 I1371 (nwayMuxOut_23n[18], inp_23d[18], nwaySelect_0n[23]);
  ND2 I1372 (nwayMuxOut_23n[19], inp_23d[19], nwaySelect_0n[23]);
  ND2 I1373 (nwayMuxOut_23n[20], inp_23d[20], nwaySelect_0n[23]);
  ND2 I1374 (nwayMuxOut_23n[21], inp_23d[21], nwaySelect_0n[23]);
  ND2 I1375 (nwayMuxOut_23n[22], inp_23d[22], nwaySelect_0n[23]);
  ND2 I1376 (nwayMuxOut_23n[23], inp_23d[23], nwaySelect_0n[23]);
  ND2 I1377 (nwayMuxOut_23n[24], inp_23d[24], nwaySelect_0n[23]);
  ND2 I1378 (nwayMuxOut_23n[25], inp_23d[25], nwaySelect_0n[23]);
  ND2 I1379 (nwayMuxOut_23n[26], inp_23d[26], nwaySelect_0n[23]);
  ND2 I1380 (nwayMuxOut_23n[27], inp_23d[27], nwaySelect_0n[23]);
  ND2 I1381 (nwayMuxOut_23n[28], inp_23d[28], nwaySelect_0n[23]);
  ND2 I1382 (nwayMuxOut_23n[29], inp_23d[29], nwaySelect_0n[23]);
  ND2 I1383 (nwayMuxOut_23n[30], inp_23d[30], nwaySelect_0n[23]);
  ND2 I1384 (nwayMuxOut_23n[31], inp_23d[31], nwaySelect_0n[23]);
  ND2 I1385 (nwayMuxOut_23n[32], inp_23d[32], nwaySelect_0n[23]);
  ND2 I1386 (nwayMuxOut_24n[0], inp_24d[0], nwaySelect_0n[24]);
  ND2 I1387 (nwayMuxOut_24n[1], inp_24d[1], nwaySelect_0n[24]);
  ND2 I1388 (nwayMuxOut_24n[2], inp_24d[2], nwaySelect_0n[24]);
  ND2 I1389 (nwayMuxOut_24n[3], inp_24d[3], nwaySelect_0n[24]);
  ND2 I1390 (nwayMuxOut_24n[4], inp_24d[4], nwaySelect_0n[24]);
  ND2 I1391 (nwayMuxOut_24n[5], inp_24d[5], nwaySelect_0n[24]);
  ND2 I1392 (nwayMuxOut_24n[6], inp_24d[6], nwaySelect_0n[24]);
  ND2 I1393 (nwayMuxOut_24n[7], inp_24d[7], nwaySelect_0n[24]);
  ND2 I1394 (nwayMuxOut_24n[8], inp_24d[8], nwaySelect_0n[24]);
  ND2 I1395 (nwayMuxOut_24n[9], inp_24d[9], nwaySelect_0n[24]);
  ND2 I1396 (nwayMuxOut_24n[10], inp_24d[10], nwaySelect_0n[24]);
  ND2 I1397 (nwayMuxOut_24n[11], inp_24d[11], nwaySelect_0n[24]);
  ND2 I1398 (nwayMuxOut_24n[12], inp_24d[12], nwaySelect_0n[24]);
  ND2 I1399 (nwayMuxOut_24n[13], inp_24d[13], nwaySelect_0n[24]);
  ND2 I1400 (nwayMuxOut_24n[14], inp_24d[14], nwaySelect_0n[24]);
  ND2 I1401 (nwayMuxOut_24n[15], inp_24d[15], nwaySelect_0n[24]);
  ND2 I1402 (nwayMuxOut_24n[16], inp_24d[16], nwaySelect_0n[24]);
  ND2 I1403 (nwayMuxOut_24n[17], inp_24d[17], nwaySelect_0n[24]);
  ND2 I1404 (nwayMuxOut_24n[18], inp_24d[18], nwaySelect_0n[24]);
  ND2 I1405 (nwayMuxOut_24n[19], inp_24d[19], nwaySelect_0n[24]);
  ND2 I1406 (nwayMuxOut_24n[20], inp_24d[20], nwaySelect_0n[24]);
  ND2 I1407 (nwayMuxOut_24n[21], inp_24d[21], nwaySelect_0n[24]);
  ND2 I1408 (nwayMuxOut_24n[22], inp_24d[22], nwaySelect_0n[24]);
  ND2 I1409 (nwayMuxOut_24n[23], inp_24d[23], nwaySelect_0n[24]);
  ND2 I1410 (nwayMuxOut_24n[24], inp_24d[24], nwaySelect_0n[24]);
  ND2 I1411 (nwayMuxOut_24n[25], inp_24d[25], nwaySelect_0n[24]);
  ND2 I1412 (nwayMuxOut_24n[26], inp_24d[26], nwaySelect_0n[24]);
  ND2 I1413 (nwayMuxOut_24n[27], inp_24d[27], nwaySelect_0n[24]);
  ND2 I1414 (nwayMuxOut_24n[28], inp_24d[28], nwaySelect_0n[24]);
  ND2 I1415 (nwayMuxOut_24n[29], inp_24d[29], nwaySelect_0n[24]);
  ND2 I1416 (nwayMuxOut_24n[30], inp_24d[30], nwaySelect_0n[24]);
  ND2 I1417 (nwayMuxOut_24n[31], inp_24d[31], nwaySelect_0n[24]);
  ND2 I1418 (nwayMuxOut_24n[32], inp_24d[32], nwaySelect_0n[24]);
  ND2 I1419 (nwayMuxOut_25n[0], inp_25d[0], nwaySelect_0n[25]);
  ND2 I1420 (nwayMuxOut_25n[1], inp_25d[1], nwaySelect_0n[25]);
  ND2 I1421 (nwayMuxOut_25n[2], inp_25d[2], nwaySelect_0n[25]);
  ND2 I1422 (nwayMuxOut_25n[3], inp_25d[3], nwaySelect_0n[25]);
  ND2 I1423 (nwayMuxOut_25n[4], inp_25d[4], nwaySelect_0n[25]);
  ND2 I1424 (nwayMuxOut_25n[5], inp_25d[5], nwaySelect_0n[25]);
  ND2 I1425 (nwayMuxOut_25n[6], inp_25d[6], nwaySelect_0n[25]);
  ND2 I1426 (nwayMuxOut_25n[7], inp_25d[7], nwaySelect_0n[25]);
  ND2 I1427 (nwayMuxOut_25n[8], inp_25d[8], nwaySelect_0n[25]);
  ND2 I1428 (nwayMuxOut_25n[9], inp_25d[9], nwaySelect_0n[25]);
  ND2 I1429 (nwayMuxOut_25n[10], inp_25d[10], nwaySelect_0n[25]);
  ND2 I1430 (nwayMuxOut_25n[11], inp_25d[11], nwaySelect_0n[25]);
  ND2 I1431 (nwayMuxOut_25n[12], inp_25d[12], nwaySelect_0n[25]);
  ND2 I1432 (nwayMuxOut_25n[13], inp_25d[13], nwaySelect_0n[25]);
  ND2 I1433 (nwayMuxOut_25n[14], inp_25d[14], nwaySelect_0n[25]);
  ND2 I1434 (nwayMuxOut_25n[15], inp_25d[15], nwaySelect_0n[25]);
  ND2 I1435 (nwayMuxOut_25n[16], inp_25d[16], nwaySelect_0n[25]);
  ND2 I1436 (nwayMuxOut_25n[17], inp_25d[17], nwaySelect_0n[25]);
  ND2 I1437 (nwayMuxOut_25n[18], inp_25d[18], nwaySelect_0n[25]);
  ND2 I1438 (nwayMuxOut_25n[19], inp_25d[19], nwaySelect_0n[25]);
  ND2 I1439 (nwayMuxOut_25n[20], inp_25d[20], nwaySelect_0n[25]);
  ND2 I1440 (nwayMuxOut_25n[21], inp_25d[21], nwaySelect_0n[25]);
  ND2 I1441 (nwayMuxOut_25n[22], inp_25d[22], nwaySelect_0n[25]);
  ND2 I1442 (nwayMuxOut_25n[23], inp_25d[23], nwaySelect_0n[25]);
  ND2 I1443 (nwayMuxOut_25n[24], inp_25d[24], nwaySelect_0n[25]);
  ND2 I1444 (nwayMuxOut_25n[25], inp_25d[25], nwaySelect_0n[25]);
  ND2 I1445 (nwayMuxOut_25n[26], inp_25d[26], nwaySelect_0n[25]);
  ND2 I1446 (nwayMuxOut_25n[27], inp_25d[27], nwaySelect_0n[25]);
  ND2 I1447 (nwayMuxOut_25n[28], inp_25d[28], nwaySelect_0n[25]);
  ND2 I1448 (nwayMuxOut_25n[29], inp_25d[29], nwaySelect_0n[25]);
  ND2 I1449 (nwayMuxOut_25n[30], inp_25d[30], nwaySelect_0n[25]);
  ND2 I1450 (nwayMuxOut_25n[31], inp_25d[31], nwaySelect_0n[25]);
  ND2 I1451 (nwayMuxOut_25n[32], inp_25d[32], nwaySelect_0n[25]);
  ND2 I1452 (nwayMuxOut_26n[0], inp_26d[0], nwaySelect_0n[26]);
  ND2 I1453 (nwayMuxOut_26n[1], inp_26d[1], nwaySelect_0n[26]);
  ND2 I1454 (nwayMuxOut_26n[2], inp_26d[2], nwaySelect_0n[26]);
  ND2 I1455 (nwayMuxOut_26n[3], inp_26d[3], nwaySelect_0n[26]);
  ND2 I1456 (nwayMuxOut_26n[4], inp_26d[4], nwaySelect_0n[26]);
  ND2 I1457 (nwayMuxOut_26n[5], inp_26d[5], nwaySelect_0n[26]);
  ND2 I1458 (nwayMuxOut_26n[6], inp_26d[6], nwaySelect_0n[26]);
  ND2 I1459 (nwayMuxOut_26n[7], inp_26d[7], nwaySelect_0n[26]);
  ND2 I1460 (nwayMuxOut_26n[8], inp_26d[8], nwaySelect_0n[26]);
  ND2 I1461 (nwayMuxOut_26n[9], inp_26d[9], nwaySelect_0n[26]);
  ND2 I1462 (nwayMuxOut_26n[10], inp_26d[10], nwaySelect_0n[26]);
  ND2 I1463 (nwayMuxOut_26n[11], inp_26d[11], nwaySelect_0n[26]);
  ND2 I1464 (nwayMuxOut_26n[12], inp_26d[12], nwaySelect_0n[26]);
  ND2 I1465 (nwayMuxOut_26n[13], inp_26d[13], nwaySelect_0n[26]);
  ND2 I1466 (nwayMuxOut_26n[14], inp_26d[14], nwaySelect_0n[26]);
  ND2 I1467 (nwayMuxOut_26n[15], inp_26d[15], nwaySelect_0n[26]);
  ND2 I1468 (nwayMuxOut_26n[16], inp_26d[16], nwaySelect_0n[26]);
  ND2 I1469 (nwayMuxOut_26n[17], inp_26d[17], nwaySelect_0n[26]);
  ND2 I1470 (nwayMuxOut_26n[18], inp_26d[18], nwaySelect_0n[26]);
  ND2 I1471 (nwayMuxOut_26n[19], inp_26d[19], nwaySelect_0n[26]);
  ND2 I1472 (nwayMuxOut_26n[20], inp_26d[20], nwaySelect_0n[26]);
  ND2 I1473 (nwayMuxOut_26n[21], inp_26d[21], nwaySelect_0n[26]);
  ND2 I1474 (nwayMuxOut_26n[22], inp_26d[22], nwaySelect_0n[26]);
  ND2 I1475 (nwayMuxOut_26n[23], inp_26d[23], nwaySelect_0n[26]);
  ND2 I1476 (nwayMuxOut_26n[24], inp_26d[24], nwaySelect_0n[26]);
  ND2 I1477 (nwayMuxOut_26n[25], inp_26d[25], nwaySelect_0n[26]);
  ND2 I1478 (nwayMuxOut_26n[26], inp_26d[26], nwaySelect_0n[26]);
  ND2 I1479 (nwayMuxOut_26n[27], inp_26d[27], nwaySelect_0n[26]);
  ND2 I1480 (nwayMuxOut_26n[28], inp_26d[28], nwaySelect_0n[26]);
  ND2 I1481 (nwayMuxOut_26n[29], inp_26d[29], nwaySelect_0n[26]);
  ND2 I1482 (nwayMuxOut_26n[30], inp_26d[30], nwaySelect_0n[26]);
  ND2 I1483 (nwayMuxOut_26n[31], inp_26d[31], nwaySelect_0n[26]);
  ND2 I1484 (nwayMuxOut_26n[32], inp_26d[32], nwaySelect_0n[26]);
  ND2 I1485 (nwayMuxOut_27n[0], inp_27d[0], nwaySelect_0n[27]);
  ND2 I1486 (nwayMuxOut_27n[1], inp_27d[1], nwaySelect_0n[27]);
  ND2 I1487 (nwayMuxOut_27n[2], inp_27d[2], nwaySelect_0n[27]);
  ND2 I1488 (nwayMuxOut_27n[3], inp_27d[3], nwaySelect_0n[27]);
  ND2 I1489 (nwayMuxOut_27n[4], inp_27d[4], nwaySelect_0n[27]);
  ND2 I1490 (nwayMuxOut_27n[5], inp_27d[5], nwaySelect_0n[27]);
  ND2 I1491 (nwayMuxOut_27n[6], inp_27d[6], nwaySelect_0n[27]);
  ND2 I1492 (nwayMuxOut_27n[7], inp_27d[7], nwaySelect_0n[27]);
  ND2 I1493 (nwayMuxOut_27n[8], inp_27d[8], nwaySelect_0n[27]);
  ND2 I1494 (nwayMuxOut_27n[9], inp_27d[9], nwaySelect_0n[27]);
  ND2 I1495 (nwayMuxOut_27n[10], inp_27d[10], nwaySelect_0n[27]);
  ND2 I1496 (nwayMuxOut_27n[11], inp_27d[11], nwaySelect_0n[27]);
  ND2 I1497 (nwayMuxOut_27n[12], inp_27d[12], nwaySelect_0n[27]);
  ND2 I1498 (nwayMuxOut_27n[13], inp_27d[13], nwaySelect_0n[27]);
  ND2 I1499 (nwayMuxOut_27n[14], inp_27d[14], nwaySelect_0n[27]);
  ND2 I1500 (nwayMuxOut_27n[15], inp_27d[15], nwaySelect_0n[27]);
  ND2 I1501 (nwayMuxOut_27n[16], inp_27d[16], nwaySelect_0n[27]);
  ND2 I1502 (nwayMuxOut_27n[17], inp_27d[17], nwaySelect_0n[27]);
  ND2 I1503 (nwayMuxOut_27n[18], inp_27d[18], nwaySelect_0n[27]);
  ND2 I1504 (nwayMuxOut_27n[19], inp_27d[19], nwaySelect_0n[27]);
  ND2 I1505 (nwayMuxOut_27n[20], inp_27d[20], nwaySelect_0n[27]);
  ND2 I1506 (nwayMuxOut_27n[21], inp_27d[21], nwaySelect_0n[27]);
  ND2 I1507 (nwayMuxOut_27n[22], inp_27d[22], nwaySelect_0n[27]);
  ND2 I1508 (nwayMuxOut_27n[23], inp_27d[23], nwaySelect_0n[27]);
  ND2 I1509 (nwayMuxOut_27n[24], inp_27d[24], nwaySelect_0n[27]);
  ND2 I1510 (nwayMuxOut_27n[25], inp_27d[25], nwaySelect_0n[27]);
  ND2 I1511 (nwayMuxOut_27n[26], inp_27d[26], nwaySelect_0n[27]);
  ND2 I1512 (nwayMuxOut_27n[27], inp_27d[27], nwaySelect_0n[27]);
  ND2 I1513 (nwayMuxOut_27n[28], inp_27d[28], nwaySelect_0n[27]);
  ND2 I1514 (nwayMuxOut_27n[29], inp_27d[29], nwaySelect_0n[27]);
  ND2 I1515 (nwayMuxOut_27n[30], inp_27d[30], nwaySelect_0n[27]);
  ND2 I1516 (nwayMuxOut_27n[31], inp_27d[31], nwaySelect_0n[27]);
  ND2 I1517 (nwayMuxOut_27n[32], inp_27d[32], nwaySelect_0n[27]);
  ND2 I1518 (nwayMuxOut_28n[0], inp_28d[0], nwaySelect_0n[28]);
  ND2 I1519 (nwayMuxOut_28n[1], inp_28d[1], nwaySelect_0n[28]);
  ND2 I1520 (nwayMuxOut_28n[2], inp_28d[2], nwaySelect_0n[28]);
  ND2 I1521 (nwayMuxOut_28n[3], inp_28d[3], nwaySelect_0n[28]);
  ND2 I1522 (nwayMuxOut_28n[4], inp_28d[4], nwaySelect_0n[28]);
  ND2 I1523 (nwayMuxOut_28n[5], inp_28d[5], nwaySelect_0n[28]);
  ND2 I1524 (nwayMuxOut_28n[6], inp_28d[6], nwaySelect_0n[28]);
  ND2 I1525 (nwayMuxOut_28n[7], inp_28d[7], nwaySelect_0n[28]);
  ND2 I1526 (nwayMuxOut_28n[8], inp_28d[8], nwaySelect_0n[28]);
  ND2 I1527 (nwayMuxOut_28n[9], inp_28d[9], nwaySelect_0n[28]);
  ND2 I1528 (nwayMuxOut_28n[10], inp_28d[10], nwaySelect_0n[28]);
  ND2 I1529 (nwayMuxOut_28n[11], inp_28d[11], nwaySelect_0n[28]);
  ND2 I1530 (nwayMuxOut_28n[12], inp_28d[12], nwaySelect_0n[28]);
  ND2 I1531 (nwayMuxOut_28n[13], inp_28d[13], nwaySelect_0n[28]);
  ND2 I1532 (nwayMuxOut_28n[14], inp_28d[14], nwaySelect_0n[28]);
  ND2 I1533 (nwayMuxOut_28n[15], inp_28d[15], nwaySelect_0n[28]);
  ND2 I1534 (nwayMuxOut_28n[16], inp_28d[16], nwaySelect_0n[28]);
  ND2 I1535 (nwayMuxOut_28n[17], inp_28d[17], nwaySelect_0n[28]);
  ND2 I1536 (nwayMuxOut_28n[18], inp_28d[18], nwaySelect_0n[28]);
  ND2 I1537 (nwayMuxOut_28n[19], inp_28d[19], nwaySelect_0n[28]);
  ND2 I1538 (nwayMuxOut_28n[20], inp_28d[20], nwaySelect_0n[28]);
  ND2 I1539 (nwayMuxOut_28n[21], inp_28d[21], nwaySelect_0n[28]);
  ND2 I1540 (nwayMuxOut_28n[22], inp_28d[22], nwaySelect_0n[28]);
  ND2 I1541 (nwayMuxOut_28n[23], inp_28d[23], nwaySelect_0n[28]);
  ND2 I1542 (nwayMuxOut_28n[24], inp_28d[24], nwaySelect_0n[28]);
  ND2 I1543 (nwayMuxOut_28n[25], inp_28d[25], nwaySelect_0n[28]);
  ND2 I1544 (nwayMuxOut_28n[26], inp_28d[26], nwaySelect_0n[28]);
  ND2 I1545 (nwayMuxOut_28n[27], inp_28d[27], nwaySelect_0n[28]);
  ND2 I1546 (nwayMuxOut_28n[28], inp_28d[28], nwaySelect_0n[28]);
  ND2 I1547 (nwayMuxOut_28n[29], inp_28d[29], nwaySelect_0n[28]);
  ND2 I1548 (nwayMuxOut_28n[30], inp_28d[30], nwaySelect_0n[28]);
  ND2 I1549 (nwayMuxOut_28n[31], inp_28d[31], nwaySelect_0n[28]);
  ND2 I1550 (nwayMuxOut_28n[32], inp_28d[32], nwaySelect_0n[28]);
  ND2 I1551 (nwayMuxOut_29n[0], inp_29d[0], nwaySelect_0n[29]);
  ND2 I1552 (nwayMuxOut_29n[1], inp_29d[1], nwaySelect_0n[29]);
  ND2 I1553 (nwayMuxOut_29n[2], inp_29d[2], nwaySelect_0n[29]);
  ND2 I1554 (nwayMuxOut_29n[3], inp_29d[3], nwaySelect_0n[29]);
  ND2 I1555 (nwayMuxOut_29n[4], inp_29d[4], nwaySelect_0n[29]);
  ND2 I1556 (nwayMuxOut_29n[5], inp_29d[5], nwaySelect_0n[29]);
  ND2 I1557 (nwayMuxOut_29n[6], inp_29d[6], nwaySelect_0n[29]);
  ND2 I1558 (nwayMuxOut_29n[7], inp_29d[7], nwaySelect_0n[29]);
  ND2 I1559 (nwayMuxOut_29n[8], inp_29d[8], nwaySelect_0n[29]);
  ND2 I1560 (nwayMuxOut_29n[9], inp_29d[9], nwaySelect_0n[29]);
  ND2 I1561 (nwayMuxOut_29n[10], inp_29d[10], nwaySelect_0n[29]);
  ND2 I1562 (nwayMuxOut_29n[11], inp_29d[11], nwaySelect_0n[29]);
  ND2 I1563 (nwayMuxOut_29n[12], inp_29d[12], nwaySelect_0n[29]);
  ND2 I1564 (nwayMuxOut_29n[13], inp_29d[13], nwaySelect_0n[29]);
  ND2 I1565 (nwayMuxOut_29n[14], inp_29d[14], nwaySelect_0n[29]);
  ND2 I1566 (nwayMuxOut_29n[15], inp_29d[15], nwaySelect_0n[29]);
  ND2 I1567 (nwayMuxOut_29n[16], inp_29d[16], nwaySelect_0n[29]);
  ND2 I1568 (nwayMuxOut_29n[17], inp_29d[17], nwaySelect_0n[29]);
  ND2 I1569 (nwayMuxOut_29n[18], inp_29d[18], nwaySelect_0n[29]);
  ND2 I1570 (nwayMuxOut_29n[19], inp_29d[19], nwaySelect_0n[29]);
  ND2 I1571 (nwayMuxOut_29n[20], inp_29d[20], nwaySelect_0n[29]);
  ND2 I1572 (nwayMuxOut_29n[21], inp_29d[21], nwaySelect_0n[29]);
  ND2 I1573 (nwayMuxOut_29n[22], inp_29d[22], nwaySelect_0n[29]);
  ND2 I1574 (nwayMuxOut_29n[23], inp_29d[23], nwaySelect_0n[29]);
  ND2 I1575 (nwayMuxOut_29n[24], inp_29d[24], nwaySelect_0n[29]);
  ND2 I1576 (nwayMuxOut_29n[25], inp_29d[25], nwaySelect_0n[29]);
  ND2 I1577 (nwayMuxOut_29n[26], inp_29d[26], nwaySelect_0n[29]);
  ND2 I1578 (nwayMuxOut_29n[27], inp_29d[27], nwaySelect_0n[29]);
  ND2 I1579 (nwayMuxOut_29n[28], inp_29d[28], nwaySelect_0n[29]);
  ND2 I1580 (nwayMuxOut_29n[29], inp_29d[29], nwaySelect_0n[29]);
  ND2 I1581 (nwayMuxOut_29n[30], inp_29d[30], nwaySelect_0n[29]);
  ND2 I1582 (nwayMuxOut_29n[31], inp_29d[31], nwaySelect_0n[29]);
  ND2 I1583 (nwayMuxOut_29n[32], inp_29d[32], nwaySelect_0n[29]);
  ND2 I1584 (nwayMuxOut_30n[0], inp_30d[0], nwaySelect_0n[30]);
  ND2 I1585 (nwayMuxOut_30n[1], inp_30d[1], nwaySelect_0n[30]);
  ND2 I1586 (nwayMuxOut_30n[2], inp_30d[2], nwaySelect_0n[30]);
  ND2 I1587 (nwayMuxOut_30n[3], inp_30d[3], nwaySelect_0n[30]);
  ND2 I1588 (nwayMuxOut_30n[4], inp_30d[4], nwaySelect_0n[30]);
  ND2 I1589 (nwayMuxOut_30n[5], inp_30d[5], nwaySelect_0n[30]);
  ND2 I1590 (nwayMuxOut_30n[6], inp_30d[6], nwaySelect_0n[30]);
  ND2 I1591 (nwayMuxOut_30n[7], inp_30d[7], nwaySelect_0n[30]);
  ND2 I1592 (nwayMuxOut_30n[8], inp_30d[8], nwaySelect_0n[30]);
  ND2 I1593 (nwayMuxOut_30n[9], inp_30d[9], nwaySelect_0n[30]);
  ND2 I1594 (nwayMuxOut_30n[10], inp_30d[10], nwaySelect_0n[30]);
  ND2 I1595 (nwayMuxOut_30n[11], inp_30d[11], nwaySelect_0n[30]);
  ND2 I1596 (nwayMuxOut_30n[12], inp_30d[12], nwaySelect_0n[30]);
  ND2 I1597 (nwayMuxOut_30n[13], inp_30d[13], nwaySelect_0n[30]);
  ND2 I1598 (nwayMuxOut_30n[14], inp_30d[14], nwaySelect_0n[30]);
  ND2 I1599 (nwayMuxOut_30n[15], inp_30d[15], nwaySelect_0n[30]);
  ND2 I1600 (nwayMuxOut_30n[16], inp_30d[16], nwaySelect_0n[30]);
  ND2 I1601 (nwayMuxOut_30n[17], inp_30d[17], nwaySelect_0n[30]);
  ND2 I1602 (nwayMuxOut_30n[18], inp_30d[18], nwaySelect_0n[30]);
  ND2 I1603 (nwayMuxOut_30n[19], inp_30d[19], nwaySelect_0n[30]);
  ND2 I1604 (nwayMuxOut_30n[20], inp_30d[20], nwaySelect_0n[30]);
  ND2 I1605 (nwayMuxOut_30n[21], inp_30d[21], nwaySelect_0n[30]);
  ND2 I1606 (nwayMuxOut_30n[22], inp_30d[22], nwaySelect_0n[30]);
  ND2 I1607 (nwayMuxOut_30n[23], inp_30d[23], nwaySelect_0n[30]);
  ND2 I1608 (nwayMuxOut_30n[24], inp_30d[24], nwaySelect_0n[30]);
  ND2 I1609 (nwayMuxOut_30n[25], inp_30d[25], nwaySelect_0n[30]);
  ND2 I1610 (nwayMuxOut_30n[26], inp_30d[26], nwaySelect_0n[30]);
  ND2 I1611 (nwayMuxOut_30n[27], inp_30d[27], nwaySelect_0n[30]);
  ND2 I1612 (nwayMuxOut_30n[28], inp_30d[28], nwaySelect_0n[30]);
  ND2 I1613 (nwayMuxOut_30n[29], inp_30d[29], nwaySelect_0n[30]);
  ND2 I1614 (nwayMuxOut_30n[30], inp_30d[30], nwaySelect_0n[30]);
  ND2 I1615 (nwayMuxOut_30n[31], inp_30d[31], nwaySelect_0n[30]);
  ND2 I1616 (nwayMuxOut_30n[32], inp_30d[32], nwaySelect_0n[30]);
  ND2 I1617 (nwayMuxOut_31n[0], inp_31d[0], nwaySelect_0n[31]);
  ND2 I1618 (nwayMuxOut_31n[1], inp_31d[1], nwaySelect_0n[31]);
  ND2 I1619 (nwayMuxOut_31n[2], inp_31d[2], nwaySelect_0n[31]);
  ND2 I1620 (nwayMuxOut_31n[3], inp_31d[3], nwaySelect_0n[31]);
  ND2 I1621 (nwayMuxOut_31n[4], inp_31d[4], nwaySelect_0n[31]);
  ND2 I1622 (nwayMuxOut_31n[5], inp_31d[5], nwaySelect_0n[31]);
  ND2 I1623 (nwayMuxOut_31n[6], inp_31d[6], nwaySelect_0n[31]);
  ND2 I1624 (nwayMuxOut_31n[7], inp_31d[7], nwaySelect_0n[31]);
  ND2 I1625 (nwayMuxOut_31n[8], inp_31d[8], nwaySelect_0n[31]);
  ND2 I1626 (nwayMuxOut_31n[9], inp_31d[9], nwaySelect_0n[31]);
  ND2 I1627 (nwayMuxOut_31n[10], inp_31d[10], nwaySelect_0n[31]);
  ND2 I1628 (nwayMuxOut_31n[11], inp_31d[11], nwaySelect_0n[31]);
  ND2 I1629 (nwayMuxOut_31n[12], inp_31d[12], nwaySelect_0n[31]);
  ND2 I1630 (nwayMuxOut_31n[13], inp_31d[13], nwaySelect_0n[31]);
  ND2 I1631 (nwayMuxOut_31n[14], inp_31d[14], nwaySelect_0n[31]);
  ND2 I1632 (nwayMuxOut_31n[15], inp_31d[15], nwaySelect_0n[31]);
  ND2 I1633 (nwayMuxOut_31n[16], inp_31d[16], nwaySelect_0n[31]);
  ND2 I1634 (nwayMuxOut_31n[17], inp_31d[17], nwaySelect_0n[31]);
  ND2 I1635 (nwayMuxOut_31n[18], inp_31d[18], nwaySelect_0n[31]);
  ND2 I1636 (nwayMuxOut_31n[19], inp_31d[19], nwaySelect_0n[31]);
  ND2 I1637 (nwayMuxOut_31n[20], inp_31d[20], nwaySelect_0n[31]);
  ND2 I1638 (nwayMuxOut_31n[21], inp_31d[21], nwaySelect_0n[31]);
  ND2 I1639 (nwayMuxOut_31n[22], inp_31d[22], nwaySelect_0n[31]);
  ND2 I1640 (nwayMuxOut_31n[23], inp_31d[23], nwaySelect_0n[31]);
  ND2 I1641 (nwayMuxOut_31n[24], inp_31d[24], nwaySelect_0n[31]);
  ND2 I1642 (nwayMuxOut_31n[25], inp_31d[25], nwaySelect_0n[31]);
  ND2 I1643 (nwayMuxOut_31n[26], inp_31d[26], nwaySelect_0n[31]);
  ND2 I1644 (nwayMuxOut_31n[27], inp_31d[27], nwaySelect_0n[31]);
  ND2 I1645 (nwayMuxOut_31n[28], inp_31d[28], nwaySelect_0n[31]);
  ND2 I1646 (nwayMuxOut_31n[29], inp_31d[29], nwaySelect_0n[31]);
  ND2 I1647 (nwayMuxOut_31n[30], inp_31d[30], nwaySelect_0n[31]);
  ND2 I1648 (nwayMuxOut_31n[31], inp_31d[31], nwaySelect_0n[31]);
  ND2 I1649 (nwayMuxOut_31n[32], inp_31d[32], nwaySelect_0n[31]);
  ND2 I1650 (nwayMuxOut_32n[0], inp_32d[0], nwaySelect_0n[32]);
  ND2 I1651 (nwayMuxOut_32n[1], inp_32d[1], nwaySelect_0n[32]);
  ND2 I1652 (nwayMuxOut_32n[2], inp_32d[2], nwaySelect_0n[32]);
  ND2 I1653 (nwayMuxOut_32n[3], inp_32d[3], nwaySelect_0n[32]);
  ND2 I1654 (nwayMuxOut_32n[4], inp_32d[4], nwaySelect_0n[32]);
  ND2 I1655 (nwayMuxOut_32n[5], inp_32d[5], nwaySelect_0n[32]);
  ND2 I1656 (nwayMuxOut_32n[6], inp_32d[6], nwaySelect_0n[32]);
  ND2 I1657 (nwayMuxOut_32n[7], inp_32d[7], nwaySelect_0n[32]);
  ND2 I1658 (nwayMuxOut_32n[8], inp_32d[8], nwaySelect_0n[32]);
  ND2 I1659 (nwayMuxOut_32n[9], inp_32d[9], nwaySelect_0n[32]);
  ND2 I1660 (nwayMuxOut_32n[10], inp_32d[10], nwaySelect_0n[32]);
  ND2 I1661 (nwayMuxOut_32n[11], inp_32d[11], nwaySelect_0n[32]);
  ND2 I1662 (nwayMuxOut_32n[12], inp_32d[12], nwaySelect_0n[32]);
  ND2 I1663 (nwayMuxOut_32n[13], inp_32d[13], nwaySelect_0n[32]);
  ND2 I1664 (nwayMuxOut_32n[14], inp_32d[14], nwaySelect_0n[32]);
  ND2 I1665 (nwayMuxOut_32n[15], inp_32d[15], nwaySelect_0n[32]);
  ND2 I1666 (nwayMuxOut_32n[16], inp_32d[16], nwaySelect_0n[32]);
  ND2 I1667 (nwayMuxOut_32n[17], inp_32d[17], nwaySelect_0n[32]);
  ND2 I1668 (nwayMuxOut_32n[18], inp_32d[18], nwaySelect_0n[32]);
  ND2 I1669 (nwayMuxOut_32n[19], inp_32d[19], nwaySelect_0n[32]);
  ND2 I1670 (nwayMuxOut_32n[20], inp_32d[20], nwaySelect_0n[32]);
  ND2 I1671 (nwayMuxOut_32n[21], inp_32d[21], nwaySelect_0n[32]);
  ND2 I1672 (nwayMuxOut_32n[22], inp_32d[22], nwaySelect_0n[32]);
  ND2 I1673 (nwayMuxOut_32n[23], inp_32d[23], nwaySelect_0n[32]);
  ND2 I1674 (nwayMuxOut_32n[24], inp_32d[24], nwaySelect_0n[32]);
  ND2 I1675 (nwayMuxOut_32n[25], inp_32d[25], nwaySelect_0n[32]);
  ND2 I1676 (nwayMuxOut_32n[26], inp_32d[26], nwaySelect_0n[32]);
  ND2 I1677 (nwayMuxOut_32n[27], inp_32d[27], nwaySelect_0n[32]);
  ND2 I1678 (nwayMuxOut_32n[28], inp_32d[28], nwaySelect_0n[32]);
  ND2 I1679 (nwayMuxOut_32n[29], inp_32d[29], nwaySelect_0n[32]);
  ND2 I1680 (nwayMuxOut_32n[30], inp_32d[30], nwaySelect_0n[32]);
  ND2 I1681 (nwayMuxOut_32n[31], inp_32d[31], nwaySelect_0n[32]);
  ND2 I1682 (nwayMuxOut_32n[32], inp_32d[32], nwaySelect_0n[32]);
  ND2 I1683 (nwayMuxOut_33n[0], inp_33d[0], nwaySelect_0n[33]);
  ND2 I1684 (nwayMuxOut_33n[1], inp_33d[1], nwaySelect_0n[33]);
  ND2 I1685 (nwayMuxOut_33n[2], inp_33d[2], nwaySelect_0n[33]);
  ND2 I1686 (nwayMuxOut_33n[3], inp_33d[3], nwaySelect_0n[33]);
  ND2 I1687 (nwayMuxOut_33n[4], inp_33d[4], nwaySelect_0n[33]);
  ND2 I1688 (nwayMuxOut_33n[5], inp_33d[5], nwaySelect_0n[33]);
  ND2 I1689 (nwayMuxOut_33n[6], inp_33d[6], nwaySelect_0n[33]);
  ND2 I1690 (nwayMuxOut_33n[7], inp_33d[7], nwaySelect_0n[33]);
  ND2 I1691 (nwayMuxOut_33n[8], inp_33d[8], nwaySelect_0n[33]);
  ND2 I1692 (nwayMuxOut_33n[9], inp_33d[9], nwaySelect_0n[33]);
  ND2 I1693 (nwayMuxOut_33n[10], inp_33d[10], nwaySelect_0n[33]);
  ND2 I1694 (nwayMuxOut_33n[11], inp_33d[11], nwaySelect_0n[33]);
  ND2 I1695 (nwayMuxOut_33n[12], inp_33d[12], nwaySelect_0n[33]);
  ND2 I1696 (nwayMuxOut_33n[13], inp_33d[13], nwaySelect_0n[33]);
  ND2 I1697 (nwayMuxOut_33n[14], inp_33d[14], nwaySelect_0n[33]);
  ND2 I1698 (nwayMuxOut_33n[15], inp_33d[15], nwaySelect_0n[33]);
  ND2 I1699 (nwayMuxOut_33n[16], inp_33d[16], nwaySelect_0n[33]);
  ND2 I1700 (nwayMuxOut_33n[17], inp_33d[17], nwaySelect_0n[33]);
  ND2 I1701 (nwayMuxOut_33n[18], inp_33d[18], nwaySelect_0n[33]);
  ND2 I1702 (nwayMuxOut_33n[19], inp_33d[19], nwaySelect_0n[33]);
  ND2 I1703 (nwayMuxOut_33n[20], inp_33d[20], nwaySelect_0n[33]);
  ND2 I1704 (nwayMuxOut_33n[21], inp_33d[21], nwaySelect_0n[33]);
  ND2 I1705 (nwayMuxOut_33n[22], inp_33d[22], nwaySelect_0n[33]);
  ND2 I1706 (nwayMuxOut_33n[23], inp_33d[23], nwaySelect_0n[33]);
  ND2 I1707 (nwayMuxOut_33n[24], inp_33d[24], nwaySelect_0n[33]);
  ND2 I1708 (nwayMuxOut_33n[25], inp_33d[25], nwaySelect_0n[33]);
  ND2 I1709 (nwayMuxOut_33n[26], inp_33d[26], nwaySelect_0n[33]);
  ND2 I1710 (nwayMuxOut_33n[27], inp_33d[27], nwaySelect_0n[33]);
  ND2 I1711 (nwayMuxOut_33n[28], inp_33d[28], nwaySelect_0n[33]);
  ND2 I1712 (nwayMuxOut_33n[29], inp_33d[29], nwaySelect_0n[33]);
  ND2 I1713 (nwayMuxOut_33n[30], inp_33d[30], nwaySelect_0n[33]);
  ND2 I1714 (nwayMuxOut_33n[31], inp_33d[31], nwaySelect_0n[33]);
  ND2 I1715 (nwayMuxOut_33n[32], inp_33d[32], nwaySelect_0n[33]);
  ND2 I1716 (nwayMuxOut_34n[0], inp_34d[0], nwaySelect_0n[34]);
  ND2 I1717 (nwayMuxOut_34n[1], inp_34d[1], nwaySelect_0n[34]);
  ND2 I1718 (nwayMuxOut_34n[2], inp_34d[2], nwaySelect_0n[34]);
  ND2 I1719 (nwayMuxOut_34n[3], inp_34d[3], nwaySelect_0n[34]);
  ND2 I1720 (nwayMuxOut_34n[4], inp_34d[4], nwaySelect_0n[34]);
  ND2 I1721 (nwayMuxOut_34n[5], inp_34d[5], nwaySelect_0n[34]);
  ND2 I1722 (nwayMuxOut_34n[6], inp_34d[6], nwaySelect_0n[34]);
  ND2 I1723 (nwayMuxOut_34n[7], inp_34d[7], nwaySelect_0n[34]);
  ND2 I1724 (nwayMuxOut_34n[8], inp_34d[8], nwaySelect_0n[34]);
  ND2 I1725 (nwayMuxOut_34n[9], inp_34d[9], nwaySelect_0n[34]);
  ND2 I1726 (nwayMuxOut_34n[10], inp_34d[10], nwaySelect_0n[34]);
  ND2 I1727 (nwayMuxOut_34n[11], inp_34d[11], nwaySelect_0n[34]);
  ND2 I1728 (nwayMuxOut_34n[12], inp_34d[12], nwaySelect_0n[34]);
  ND2 I1729 (nwayMuxOut_34n[13], inp_34d[13], nwaySelect_0n[34]);
  ND2 I1730 (nwayMuxOut_34n[14], inp_34d[14], nwaySelect_0n[34]);
  ND2 I1731 (nwayMuxOut_34n[15], inp_34d[15], nwaySelect_0n[34]);
  ND2 I1732 (nwayMuxOut_34n[16], inp_34d[16], nwaySelect_0n[34]);
  ND2 I1733 (nwayMuxOut_34n[17], inp_34d[17], nwaySelect_0n[34]);
  ND2 I1734 (nwayMuxOut_34n[18], inp_34d[18], nwaySelect_0n[34]);
  ND2 I1735 (nwayMuxOut_34n[19], inp_34d[19], nwaySelect_0n[34]);
  ND2 I1736 (nwayMuxOut_34n[20], inp_34d[20], nwaySelect_0n[34]);
  ND2 I1737 (nwayMuxOut_34n[21], inp_34d[21], nwaySelect_0n[34]);
  ND2 I1738 (nwayMuxOut_34n[22], inp_34d[22], nwaySelect_0n[34]);
  ND2 I1739 (nwayMuxOut_34n[23], inp_34d[23], nwaySelect_0n[34]);
  ND2 I1740 (nwayMuxOut_34n[24], inp_34d[24], nwaySelect_0n[34]);
  ND2 I1741 (nwayMuxOut_34n[25], inp_34d[25], nwaySelect_0n[34]);
  ND2 I1742 (nwayMuxOut_34n[26], inp_34d[26], nwaySelect_0n[34]);
  ND2 I1743 (nwayMuxOut_34n[27], inp_34d[27], nwaySelect_0n[34]);
  ND2 I1744 (nwayMuxOut_34n[28], inp_34d[28], nwaySelect_0n[34]);
  ND2 I1745 (nwayMuxOut_34n[29], inp_34d[29], nwaySelect_0n[34]);
  ND2 I1746 (nwayMuxOut_34n[30], inp_34d[30], nwaySelect_0n[34]);
  ND2 I1747 (nwayMuxOut_34n[31], inp_34d[31], nwaySelect_0n[34]);
  ND2 I1748 (nwayMuxOut_34n[32], inp_34d[32], nwaySelect_0n[34]);
  ND2 I1749 (nwayMuxOut_35n[0], inp_35d[0], nwaySelect_0n[35]);
  ND2 I1750 (nwayMuxOut_35n[1], inp_35d[1], nwaySelect_0n[35]);
  ND2 I1751 (nwayMuxOut_35n[2], inp_35d[2], nwaySelect_0n[35]);
  ND2 I1752 (nwayMuxOut_35n[3], inp_35d[3], nwaySelect_0n[35]);
  ND2 I1753 (nwayMuxOut_35n[4], inp_35d[4], nwaySelect_0n[35]);
  ND2 I1754 (nwayMuxOut_35n[5], inp_35d[5], nwaySelect_0n[35]);
  ND2 I1755 (nwayMuxOut_35n[6], inp_35d[6], nwaySelect_0n[35]);
  ND2 I1756 (nwayMuxOut_35n[7], inp_35d[7], nwaySelect_0n[35]);
  ND2 I1757 (nwayMuxOut_35n[8], inp_35d[8], nwaySelect_0n[35]);
  ND2 I1758 (nwayMuxOut_35n[9], inp_35d[9], nwaySelect_0n[35]);
  ND2 I1759 (nwayMuxOut_35n[10], inp_35d[10], nwaySelect_0n[35]);
  ND2 I1760 (nwayMuxOut_35n[11], inp_35d[11], nwaySelect_0n[35]);
  ND2 I1761 (nwayMuxOut_35n[12], inp_35d[12], nwaySelect_0n[35]);
  ND2 I1762 (nwayMuxOut_35n[13], inp_35d[13], nwaySelect_0n[35]);
  ND2 I1763 (nwayMuxOut_35n[14], inp_35d[14], nwaySelect_0n[35]);
  ND2 I1764 (nwayMuxOut_35n[15], inp_35d[15], nwaySelect_0n[35]);
  ND2 I1765 (nwayMuxOut_35n[16], inp_35d[16], nwaySelect_0n[35]);
  ND2 I1766 (nwayMuxOut_35n[17], inp_35d[17], nwaySelect_0n[35]);
  ND2 I1767 (nwayMuxOut_35n[18], inp_35d[18], nwaySelect_0n[35]);
  ND2 I1768 (nwayMuxOut_35n[19], inp_35d[19], nwaySelect_0n[35]);
  ND2 I1769 (nwayMuxOut_35n[20], inp_35d[20], nwaySelect_0n[35]);
  ND2 I1770 (nwayMuxOut_35n[21], inp_35d[21], nwaySelect_0n[35]);
  ND2 I1771 (nwayMuxOut_35n[22], inp_35d[22], nwaySelect_0n[35]);
  ND2 I1772 (nwayMuxOut_35n[23], inp_35d[23], nwaySelect_0n[35]);
  ND2 I1773 (nwayMuxOut_35n[24], inp_35d[24], nwaySelect_0n[35]);
  ND2 I1774 (nwayMuxOut_35n[25], inp_35d[25], nwaySelect_0n[35]);
  ND2 I1775 (nwayMuxOut_35n[26], inp_35d[26], nwaySelect_0n[35]);
  ND2 I1776 (nwayMuxOut_35n[27], inp_35d[27], nwaySelect_0n[35]);
  ND2 I1777 (nwayMuxOut_35n[28], inp_35d[28], nwaySelect_0n[35]);
  ND2 I1778 (nwayMuxOut_35n[29], inp_35d[29], nwaySelect_0n[35]);
  ND2 I1779 (nwayMuxOut_35n[30], inp_35d[30], nwaySelect_0n[35]);
  ND2 I1780 (nwayMuxOut_35n[31], inp_35d[31], nwaySelect_0n[35]);
  ND2 I1781 (nwayMuxOut_35n[32], inp_35d[32], nwaySelect_0n[35]);
  ND2 I1782 (nwayMuxOut_36n[0], inp_36d[0], nwaySelect_0n[36]);
  ND2 I1783 (nwayMuxOut_36n[1], inp_36d[1], nwaySelect_0n[36]);
  ND2 I1784 (nwayMuxOut_36n[2], inp_36d[2], nwaySelect_0n[36]);
  ND2 I1785 (nwayMuxOut_36n[3], inp_36d[3], nwaySelect_0n[36]);
  ND2 I1786 (nwayMuxOut_36n[4], inp_36d[4], nwaySelect_0n[36]);
  ND2 I1787 (nwayMuxOut_36n[5], inp_36d[5], nwaySelect_0n[36]);
  ND2 I1788 (nwayMuxOut_36n[6], inp_36d[6], nwaySelect_0n[36]);
  ND2 I1789 (nwayMuxOut_36n[7], inp_36d[7], nwaySelect_0n[36]);
  ND2 I1790 (nwayMuxOut_36n[8], inp_36d[8], nwaySelect_0n[36]);
  ND2 I1791 (nwayMuxOut_36n[9], inp_36d[9], nwaySelect_0n[36]);
  ND2 I1792 (nwayMuxOut_36n[10], inp_36d[10], nwaySelect_0n[36]);
  ND2 I1793 (nwayMuxOut_36n[11], inp_36d[11], nwaySelect_0n[36]);
  ND2 I1794 (nwayMuxOut_36n[12], inp_36d[12], nwaySelect_0n[36]);
  ND2 I1795 (nwayMuxOut_36n[13], inp_36d[13], nwaySelect_0n[36]);
  ND2 I1796 (nwayMuxOut_36n[14], inp_36d[14], nwaySelect_0n[36]);
  ND2 I1797 (nwayMuxOut_36n[15], inp_36d[15], nwaySelect_0n[36]);
  ND2 I1798 (nwayMuxOut_36n[16], inp_36d[16], nwaySelect_0n[36]);
  ND2 I1799 (nwayMuxOut_36n[17], inp_36d[17], nwaySelect_0n[36]);
  ND2 I1800 (nwayMuxOut_36n[18], inp_36d[18], nwaySelect_0n[36]);
  ND2 I1801 (nwayMuxOut_36n[19], inp_36d[19], nwaySelect_0n[36]);
  ND2 I1802 (nwayMuxOut_36n[20], inp_36d[20], nwaySelect_0n[36]);
  ND2 I1803 (nwayMuxOut_36n[21], inp_36d[21], nwaySelect_0n[36]);
  ND2 I1804 (nwayMuxOut_36n[22], inp_36d[22], nwaySelect_0n[36]);
  ND2 I1805 (nwayMuxOut_36n[23], inp_36d[23], nwaySelect_0n[36]);
  ND2 I1806 (nwayMuxOut_36n[24], inp_36d[24], nwaySelect_0n[36]);
  ND2 I1807 (nwayMuxOut_36n[25], inp_36d[25], nwaySelect_0n[36]);
  ND2 I1808 (nwayMuxOut_36n[26], inp_36d[26], nwaySelect_0n[36]);
  ND2 I1809 (nwayMuxOut_36n[27], inp_36d[27], nwaySelect_0n[36]);
  ND2 I1810 (nwayMuxOut_36n[28], inp_36d[28], nwaySelect_0n[36]);
  ND2 I1811 (nwayMuxOut_36n[29], inp_36d[29], nwaySelect_0n[36]);
  ND2 I1812 (nwayMuxOut_36n[30], inp_36d[30], nwaySelect_0n[36]);
  ND2 I1813 (nwayMuxOut_36n[31], inp_36d[31], nwaySelect_0n[36]);
  ND2 I1814 (nwayMuxOut_36n[32], inp_36d[32], nwaySelect_0n[36]);
  ND2 I1815 (nwayMuxOut_37n[0], inp_37d[0], nwaySelect_0n[37]);
  ND2 I1816 (nwayMuxOut_37n[1], inp_37d[1], nwaySelect_0n[37]);
  ND2 I1817 (nwayMuxOut_37n[2], inp_37d[2], nwaySelect_0n[37]);
  ND2 I1818 (nwayMuxOut_37n[3], inp_37d[3], nwaySelect_0n[37]);
  ND2 I1819 (nwayMuxOut_37n[4], inp_37d[4], nwaySelect_0n[37]);
  ND2 I1820 (nwayMuxOut_37n[5], inp_37d[5], nwaySelect_0n[37]);
  ND2 I1821 (nwayMuxOut_37n[6], inp_37d[6], nwaySelect_0n[37]);
  ND2 I1822 (nwayMuxOut_37n[7], inp_37d[7], nwaySelect_0n[37]);
  ND2 I1823 (nwayMuxOut_37n[8], inp_37d[8], nwaySelect_0n[37]);
  ND2 I1824 (nwayMuxOut_37n[9], inp_37d[9], nwaySelect_0n[37]);
  ND2 I1825 (nwayMuxOut_37n[10], inp_37d[10], nwaySelect_0n[37]);
  ND2 I1826 (nwayMuxOut_37n[11], inp_37d[11], nwaySelect_0n[37]);
  ND2 I1827 (nwayMuxOut_37n[12], inp_37d[12], nwaySelect_0n[37]);
  ND2 I1828 (nwayMuxOut_37n[13], inp_37d[13], nwaySelect_0n[37]);
  ND2 I1829 (nwayMuxOut_37n[14], inp_37d[14], nwaySelect_0n[37]);
  ND2 I1830 (nwayMuxOut_37n[15], inp_37d[15], nwaySelect_0n[37]);
  ND2 I1831 (nwayMuxOut_37n[16], inp_37d[16], nwaySelect_0n[37]);
  ND2 I1832 (nwayMuxOut_37n[17], inp_37d[17], nwaySelect_0n[37]);
  ND2 I1833 (nwayMuxOut_37n[18], inp_37d[18], nwaySelect_0n[37]);
  ND2 I1834 (nwayMuxOut_37n[19], inp_37d[19], nwaySelect_0n[37]);
  ND2 I1835 (nwayMuxOut_37n[20], inp_37d[20], nwaySelect_0n[37]);
  ND2 I1836 (nwayMuxOut_37n[21], inp_37d[21], nwaySelect_0n[37]);
  ND2 I1837 (nwayMuxOut_37n[22], inp_37d[22], nwaySelect_0n[37]);
  ND2 I1838 (nwayMuxOut_37n[23], inp_37d[23], nwaySelect_0n[37]);
  ND2 I1839 (nwayMuxOut_37n[24], inp_37d[24], nwaySelect_0n[37]);
  ND2 I1840 (nwayMuxOut_37n[25], inp_37d[25], nwaySelect_0n[37]);
  ND2 I1841 (nwayMuxOut_37n[26], inp_37d[26], nwaySelect_0n[37]);
  ND2 I1842 (nwayMuxOut_37n[27], inp_37d[27], nwaySelect_0n[37]);
  ND2 I1843 (nwayMuxOut_37n[28], inp_37d[28], nwaySelect_0n[37]);
  ND2 I1844 (nwayMuxOut_37n[29], inp_37d[29], nwaySelect_0n[37]);
  ND2 I1845 (nwayMuxOut_37n[30], inp_37d[30], nwaySelect_0n[37]);
  ND2 I1846 (nwayMuxOut_37n[31], inp_37d[31], nwaySelect_0n[37]);
  ND2 I1847 (nwayMuxOut_37n[32], inp_37d[32], nwaySelect_0n[37]);
  ND2 I1848 (nwayMuxOut_38n[0], inp_38d[0], nwaySelect_0n[38]);
  ND2 I1849 (nwayMuxOut_38n[1], inp_38d[1], nwaySelect_0n[38]);
  ND2 I1850 (nwayMuxOut_38n[2], inp_38d[2], nwaySelect_0n[38]);
  ND2 I1851 (nwayMuxOut_38n[3], inp_38d[3], nwaySelect_0n[38]);
  ND2 I1852 (nwayMuxOut_38n[4], inp_38d[4], nwaySelect_0n[38]);
  ND2 I1853 (nwayMuxOut_38n[5], inp_38d[5], nwaySelect_0n[38]);
  ND2 I1854 (nwayMuxOut_38n[6], inp_38d[6], nwaySelect_0n[38]);
  ND2 I1855 (nwayMuxOut_38n[7], inp_38d[7], nwaySelect_0n[38]);
  ND2 I1856 (nwayMuxOut_38n[8], inp_38d[8], nwaySelect_0n[38]);
  ND2 I1857 (nwayMuxOut_38n[9], inp_38d[9], nwaySelect_0n[38]);
  ND2 I1858 (nwayMuxOut_38n[10], inp_38d[10], nwaySelect_0n[38]);
  ND2 I1859 (nwayMuxOut_38n[11], inp_38d[11], nwaySelect_0n[38]);
  ND2 I1860 (nwayMuxOut_38n[12], inp_38d[12], nwaySelect_0n[38]);
  ND2 I1861 (nwayMuxOut_38n[13], inp_38d[13], nwaySelect_0n[38]);
  ND2 I1862 (nwayMuxOut_38n[14], inp_38d[14], nwaySelect_0n[38]);
  ND2 I1863 (nwayMuxOut_38n[15], inp_38d[15], nwaySelect_0n[38]);
  ND2 I1864 (nwayMuxOut_38n[16], inp_38d[16], nwaySelect_0n[38]);
  ND2 I1865 (nwayMuxOut_38n[17], inp_38d[17], nwaySelect_0n[38]);
  ND2 I1866 (nwayMuxOut_38n[18], inp_38d[18], nwaySelect_0n[38]);
  ND2 I1867 (nwayMuxOut_38n[19], inp_38d[19], nwaySelect_0n[38]);
  ND2 I1868 (nwayMuxOut_38n[20], inp_38d[20], nwaySelect_0n[38]);
  ND2 I1869 (nwayMuxOut_38n[21], inp_38d[21], nwaySelect_0n[38]);
  ND2 I1870 (nwayMuxOut_38n[22], inp_38d[22], nwaySelect_0n[38]);
  ND2 I1871 (nwayMuxOut_38n[23], inp_38d[23], nwaySelect_0n[38]);
  ND2 I1872 (nwayMuxOut_38n[24], inp_38d[24], nwaySelect_0n[38]);
  ND2 I1873 (nwayMuxOut_38n[25], inp_38d[25], nwaySelect_0n[38]);
  ND2 I1874 (nwayMuxOut_38n[26], inp_38d[26], nwaySelect_0n[38]);
  ND2 I1875 (nwayMuxOut_38n[27], inp_38d[27], nwaySelect_0n[38]);
  ND2 I1876 (nwayMuxOut_38n[28], inp_38d[28], nwaySelect_0n[38]);
  ND2 I1877 (nwayMuxOut_38n[29], inp_38d[29], nwaySelect_0n[38]);
  ND2 I1878 (nwayMuxOut_38n[30], inp_38d[30], nwaySelect_0n[38]);
  ND2 I1879 (nwayMuxOut_38n[31], inp_38d[31], nwaySelect_0n[38]);
  ND2 I1880 (nwayMuxOut_38n[32], inp_38d[32], nwaySelect_0n[38]);
  ND2 I1881 (nwayMuxOut_39n[0], inp_39d[0], nwaySelect_0n[39]);
  ND2 I1882 (nwayMuxOut_39n[1], inp_39d[1], nwaySelect_0n[39]);
  ND2 I1883 (nwayMuxOut_39n[2], inp_39d[2], nwaySelect_0n[39]);
  ND2 I1884 (nwayMuxOut_39n[3], inp_39d[3], nwaySelect_0n[39]);
  ND2 I1885 (nwayMuxOut_39n[4], inp_39d[4], nwaySelect_0n[39]);
  ND2 I1886 (nwayMuxOut_39n[5], inp_39d[5], nwaySelect_0n[39]);
  ND2 I1887 (nwayMuxOut_39n[6], inp_39d[6], nwaySelect_0n[39]);
  ND2 I1888 (nwayMuxOut_39n[7], inp_39d[7], nwaySelect_0n[39]);
  ND2 I1889 (nwayMuxOut_39n[8], inp_39d[8], nwaySelect_0n[39]);
  ND2 I1890 (nwayMuxOut_39n[9], inp_39d[9], nwaySelect_0n[39]);
  ND2 I1891 (nwayMuxOut_39n[10], inp_39d[10], nwaySelect_0n[39]);
  ND2 I1892 (nwayMuxOut_39n[11], inp_39d[11], nwaySelect_0n[39]);
  ND2 I1893 (nwayMuxOut_39n[12], inp_39d[12], nwaySelect_0n[39]);
  ND2 I1894 (nwayMuxOut_39n[13], inp_39d[13], nwaySelect_0n[39]);
  ND2 I1895 (nwayMuxOut_39n[14], inp_39d[14], nwaySelect_0n[39]);
  ND2 I1896 (nwayMuxOut_39n[15], inp_39d[15], nwaySelect_0n[39]);
  ND2 I1897 (nwayMuxOut_39n[16], inp_39d[16], nwaySelect_0n[39]);
  ND2 I1898 (nwayMuxOut_39n[17], inp_39d[17], nwaySelect_0n[39]);
  ND2 I1899 (nwayMuxOut_39n[18], inp_39d[18], nwaySelect_0n[39]);
  ND2 I1900 (nwayMuxOut_39n[19], inp_39d[19], nwaySelect_0n[39]);
  ND2 I1901 (nwayMuxOut_39n[20], inp_39d[20], nwaySelect_0n[39]);
  ND2 I1902 (nwayMuxOut_39n[21], inp_39d[21], nwaySelect_0n[39]);
  ND2 I1903 (nwayMuxOut_39n[22], inp_39d[22], nwaySelect_0n[39]);
  ND2 I1904 (nwayMuxOut_39n[23], inp_39d[23], nwaySelect_0n[39]);
  ND2 I1905 (nwayMuxOut_39n[24], inp_39d[24], nwaySelect_0n[39]);
  ND2 I1906 (nwayMuxOut_39n[25], inp_39d[25], nwaySelect_0n[39]);
  ND2 I1907 (nwayMuxOut_39n[26], inp_39d[26], nwaySelect_0n[39]);
  ND2 I1908 (nwayMuxOut_39n[27], inp_39d[27], nwaySelect_0n[39]);
  ND2 I1909 (nwayMuxOut_39n[28], inp_39d[28], nwaySelect_0n[39]);
  ND2 I1910 (nwayMuxOut_39n[29], inp_39d[29], nwaySelect_0n[39]);
  ND2 I1911 (nwayMuxOut_39n[30], inp_39d[30], nwaySelect_0n[39]);
  ND2 I1912 (nwayMuxOut_39n[31], inp_39d[31], nwaySelect_0n[39]);
  ND2 I1913 (nwayMuxOut_39n[32], inp_39d[32], nwaySelect_0n[39]);
  ND2 I1914 (nwayMuxOut_40n[0], inp_40d[0], nwaySelect_0n[40]);
  ND2 I1915 (nwayMuxOut_40n[1], inp_40d[1], nwaySelect_0n[40]);
  ND2 I1916 (nwayMuxOut_40n[2], inp_40d[2], nwaySelect_0n[40]);
  ND2 I1917 (nwayMuxOut_40n[3], inp_40d[3], nwaySelect_0n[40]);
  ND2 I1918 (nwayMuxOut_40n[4], inp_40d[4], nwaySelect_0n[40]);
  ND2 I1919 (nwayMuxOut_40n[5], inp_40d[5], nwaySelect_0n[40]);
  ND2 I1920 (nwayMuxOut_40n[6], inp_40d[6], nwaySelect_0n[40]);
  ND2 I1921 (nwayMuxOut_40n[7], inp_40d[7], nwaySelect_0n[40]);
  ND2 I1922 (nwayMuxOut_40n[8], inp_40d[8], nwaySelect_0n[40]);
  ND2 I1923 (nwayMuxOut_40n[9], inp_40d[9], nwaySelect_0n[40]);
  ND2 I1924 (nwayMuxOut_40n[10], inp_40d[10], nwaySelect_0n[40]);
  ND2 I1925 (nwayMuxOut_40n[11], inp_40d[11], nwaySelect_0n[40]);
  ND2 I1926 (nwayMuxOut_40n[12], inp_40d[12], nwaySelect_0n[40]);
  ND2 I1927 (nwayMuxOut_40n[13], inp_40d[13], nwaySelect_0n[40]);
  ND2 I1928 (nwayMuxOut_40n[14], inp_40d[14], nwaySelect_0n[40]);
  ND2 I1929 (nwayMuxOut_40n[15], inp_40d[15], nwaySelect_0n[40]);
  ND2 I1930 (nwayMuxOut_40n[16], inp_40d[16], nwaySelect_0n[40]);
  ND2 I1931 (nwayMuxOut_40n[17], inp_40d[17], nwaySelect_0n[40]);
  ND2 I1932 (nwayMuxOut_40n[18], inp_40d[18], nwaySelect_0n[40]);
  ND2 I1933 (nwayMuxOut_40n[19], inp_40d[19], nwaySelect_0n[40]);
  ND2 I1934 (nwayMuxOut_40n[20], inp_40d[20], nwaySelect_0n[40]);
  ND2 I1935 (nwayMuxOut_40n[21], inp_40d[21], nwaySelect_0n[40]);
  ND2 I1936 (nwayMuxOut_40n[22], inp_40d[22], nwaySelect_0n[40]);
  ND2 I1937 (nwayMuxOut_40n[23], inp_40d[23], nwaySelect_0n[40]);
  ND2 I1938 (nwayMuxOut_40n[24], inp_40d[24], nwaySelect_0n[40]);
  ND2 I1939 (nwayMuxOut_40n[25], inp_40d[25], nwaySelect_0n[40]);
  ND2 I1940 (nwayMuxOut_40n[26], inp_40d[26], nwaySelect_0n[40]);
  ND2 I1941 (nwayMuxOut_40n[27], inp_40d[27], nwaySelect_0n[40]);
  ND2 I1942 (nwayMuxOut_40n[28], inp_40d[28], nwaySelect_0n[40]);
  ND2 I1943 (nwayMuxOut_40n[29], inp_40d[29], nwaySelect_0n[40]);
  ND2 I1944 (nwayMuxOut_40n[30], inp_40d[30], nwaySelect_0n[40]);
  ND2 I1945 (nwayMuxOut_40n[31], inp_40d[31], nwaySelect_0n[40]);
  ND2 I1946 (nwayMuxOut_40n[32], inp_40d[32], nwaySelect_0n[40]);
  ND2 I1947 (nwayMuxOut_41n[0], inp_41d[0], nwaySelect_0n[41]);
  ND2 I1948 (nwayMuxOut_41n[1], inp_41d[1], nwaySelect_0n[41]);
  ND2 I1949 (nwayMuxOut_41n[2], inp_41d[2], nwaySelect_0n[41]);
  ND2 I1950 (nwayMuxOut_41n[3], inp_41d[3], nwaySelect_0n[41]);
  ND2 I1951 (nwayMuxOut_41n[4], inp_41d[4], nwaySelect_0n[41]);
  ND2 I1952 (nwayMuxOut_41n[5], inp_41d[5], nwaySelect_0n[41]);
  ND2 I1953 (nwayMuxOut_41n[6], inp_41d[6], nwaySelect_0n[41]);
  ND2 I1954 (nwayMuxOut_41n[7], inp_41d[7], nwaySelect_0n[41]);
  ND2 I1955 (nwayMuxOut_41n[8], inp_41d[8], nwaySelect_0n[41]);
  ND2 I1956 (nwayMuxOut_41n[9], inp_41d[9], nwaySelect_0n[41]);
  ND2 I1957 (nwayMuxOut_41n[10], inp_41d[10], nwaySelect_0n[41]);
  ND2 I1958 (nwayMuxOut_41n[11], inp_41d[11], nwaySelect_0n[41]);
  ND2 I1959 (nwayMuxOut_41n[12], inp_41d[12], nwaySelect_0n[41]);
  ND2 I1960 (nwayMuxOut_41n[13], inp_41d[13], nwaySelect_0n[41]);
  ND2 I1961 (nwayMuxOut_41n[14], inp_41d[14], nwaySelect_0n[41]);
  ND2 I1962 (nwayMuxOut_41n[15], inp_41d[15], nwaySelect_0n[41]);
  ND2 I1963 (nwayMuxOut_41n[16], inp_41d[16], nwaySelect_0n[41]);
  ND2 I1964 (nwayMuxOut_41n[17], inp_41d[17], nwaySelect_0n[41]);
  ND2 I1965 (nwayMuxOut_41n[18], inp_41d[18], nwaySelect_0n[41]);
  ND2 I1966 (nwayMuxOut_41n[19], inp_41d[19], nwaySelect_0n[41]);
  ND2 I1967 (nwayMuxOut_41n[20], inp_41d[20], nwaySelect_0n[41]);
  ND2 I1968 (nwayMuxOut_41n[21], inp_41d[21], nwaySelect_0n[41]);
  ND2 I1969 (nwayMuxOut_41n[22], inp_41d[22], nwaySelect_0n[41]);
  ND2 I1970 (nwayMuxOut_41n[23], inp_41d[23], nwaySelect_0n[41]);
  ND2 I1971 (nwayMuxOut_41n[24], inp_41d[24], nwaySelect_0n[41]);
  ND2 I1972 (nwayMuxOut_41n[25], inp_41d[25], nwaySelect_0n[41]);
  ND2 I1973 (nwayMuxOut_41n[26], inp_41d[26], nwaySelect_0n[41]);
  ND2 I1974 (nwayMuxOut_41n[27], inp_41d[27], nwaySelect_0n[41]);
  ND2 I1975 (nwayMuxOut_41n[28], inp_41d[28], nwaySelect_0n[41]);
  ND2 I1976 (nwayMuxOut_41n[29], inp_41d[29], nwaySelect_0n[41]);
  ND2 I1977 (nwayMuxOut_41n[30], inp_41d[30], nwaySelect_0n[41]);
  ND2 I1978 (nwayMuxOut_41n[31], inp_41d[31], nwaySelect_0n[41]);
  ND2 I1979 (nwayMuxOut_41n[32], inp_41d[32], nwaySelect_0n[41]);
  ND2 I1980 (nwayMuxOut_42n[0], inp_42d[0], nwaySelect_0n[42]);
  ND2 I1981 (nwayMuxOut_42n[1], inp_42d[1], nwaySelect_0n[42]);
  ND2 I1982 (nwayMuxOut_42n[2], inp_42d[2], nwaySelect_0n[42]);
  ND2 I1983 (nwayMuxOut_42n[3], inp_42d[3], nwaySelect_0n[42]);
  ND2 I1984 (nwayMuxOut_42n[4], inp_42d[4], nwaySelect_0n[42]);
  ND2 I1985 (nwayMuxOut_42n[5], inp_42d[5], nwaySelect_0n[42]);
  ND2 I1986 (nwayMuxOut_42n[6], inp_42d[6], nwaySelect_0n[42]);
  ND2 I1987 (nwayMuxOut_42n[7], inp_42d[7], nwaySelect_0n[42]);
  ND2 I1988 (nwayMuxOut_42n[8], inp_42d[8], nwaySelect_0n[42]);
  ND2 I1989 (nwayMuxOut_42n[9], inp_42d[9], nwaySelect_0n[42]);
  ND2 I1990 (nwayMuxOut_42n[10], inp_42d[10], nwaySelect_0n[42]);
  ND2 I1991 (nwayMuxOut_42n[11], inp_42d[11], nwaySelect_0n[42]);
  ND2 I1992 (nwayMuxOut_42n[12], inp_42d[12], nwaySelect_0n[42]);
  ND2 I1993 (nwayMuxOut_42n[13], inp_42d[13], nwaySelect_0n[42]);
  ND2 I1994 (nwayMuxOut_42n[14], inp_42d[14], nwaySelect_0n[42]);
  ND2 I1995 (nwayMuxOut_42n[15], inp_42d[15], nwaySelect_0n[42]);
  ND2 I1996 (nwayMuxOut_42n[16], inp_42d[16], nwaySelect_0n[42]);
  ND2 I1997 (nwayMuxOut_42n[17], inp_42d[17], nwaySelect_0n[42]);
  ND2 I1998 (nwayMuxOut_42n[18], inp_42d[18], nwaySelect_0n[42]);
  ND2 I1999 (nwayMuxOut_42n[19], inp_42d[19], nwaySelect_0n[42]);
  ND2 I2000 (nwayMuxOut_42n[20], inp_42d[20], nwaySelect_0n[42]);
  ND2 I2001 (nwayMuxOut_42n[21], inp_42d[21], nwaySelect_0n[42]);
  ND2 I2002 (nwayMuxOut_42n[22], inp_42d[22], nwaySelect_0n[42]);
  ND2 I2003 (nwayMuxOut_42n[23], inp_42d[23], nwaySelect_0n[42]);
  ND2 I2004 (nwayMuxOut_42n[24], inp_42d[24], nwaySelect_0n[42]);
  ND2 I2005 (nwayMuxOut_42n[25], inp_42d[25], nwaySelect_0n[42]);
  ND2 I2006 (nwayMuxOut_42n[26], inp_42d[26], nwaySelect_0n[42]);
  ND2 I2007 (nwayMuxOut_42n[27], inp_42d[27], nwaySelect_0n[42]);
  ND2 I2008 (nwayMuxOut_42n[28], inp_42d[28], nwaySelect_0n[42]);
  ND2 I2009 (nwayMuxOut_42n[29], inp_42d[29], nwaySelect_0n[42]);
  ND2 I2010 (nwayMuxOut_42n[30], inp_42d[30], nwaySelect_0n[42]);
  ND2 I2011 (nwayMuxOut_42n[31], inp_42d[31], nwaySelect_0n[42]);
  ND2 I2012 (nwayMuxOut_42n[32], inp_42d[32], nwaySelect_0n[42]);
  ND2 I2013 (nwayMuxOut_43n[0], inp_43d[0], nwaySelect_0n[43]);
  ND2 I2014 (nwayMuxOut_43n[1], inp_43d[1], nwaySelect_0n[43]);
  ND2 I2015 (nwayMuxOut_43n[2], inp_43d[2], nwaySelect_0n[43]);
  ND2 I2016 (nwayMuxOut_43n[3], inp_43d[3], nwaySelect_0n[43]);
  ND2 I2017 (nwayMuxOut_43n[4], inp_43d[4], nwaySelect_0n[43]);
  ND2 I2018 (nwayMuxOut_43n[5], inp_43d[5], nwaySelect_0n[43]);
  ND2 I2019 (nwayMuxOut_43n[6], inp_43d[6], nwaySelect_0n[43]);
  ND2 I2020 (nwayMuxOut_43n[7], inp_43d[7], nwaySelect_0n[43]);
  ND2 I2021 (nwayMuxOut_43n[8], inp_43d[8], nwaySelect_0n[43]);
  ND2 I2022 (nwayMuxOut_43n[9], inp_43d[9], nwaySelect_0n[43]);
  ND2 I2023 (nwayMuxOut_43n[10], inp_43d[10], nwaySelect_0n[43]);
  ND2 I2024 (nwayMuxOut_43n[11], inp_43d[11], nwaySelect_0n[43]);
  ND2 I2025 (nwayMuxOut_43n[12], inp_43d[12], nwaySelect_0n[43]);
  ND2 I2026 (nwayMuxOut_43n[13], inp_43d[13], nwaySelect_0n[43]);
  ND2 I2027 (nwayMuxOut_43n[14], inp_43d[14], nwaySelect_0n[43]);
  ND2 I2028 (nwayMuxOut_43n[15], inp_43d[15], nwaySelect_0n[43]);
  ND2 I2029 (nwayMuxOut_43n[16], inp_43d[16], nwaySelect_0n[43]);
  ND2 I2030 (nwayMuxOut_43n[17], inp_43d[17], nwaySelect_0n[43]);
  ND2 I2031 (nwayMuxOut_43n[18], inp_43d[18], nwaySelect_0n[43]);
  ND2 I2032 (nwayMuxOut_43n[19], inp_43d[19], nwaySelect_0n[43]);
  ND2 I2033 (nwayMuxOut_43n[20], inp_43d[20], nwaySelect_0n[43]);
  ND2 I2034 (nwayMuxOut_43n[21], inp_43d[21], nwaySelect_0n[43]);
  ND2 I2035 (nwayMuxOut_43n[22], inp_43d[22], nwaySelect_0n[43]);
  ND2 I2036 (nwayMuxOut_43n[23], inp_43d[23], nwaySelect_0n[43]);
  ND2 I2037 (nwayMuxOut_43n[24], inp_43d[24], nwaySelect_0n[43]);
  ND2 I2038 (nwayMuxOut_43n[25], inp_43d[25], nwaySelect_0n[43]);
  ND2 I2039 (nwayMuxOut_43n[26], inp_43d[26], nwaySelect_0n[43]);
  ND2 I2040 (nwayMuxOut_43n[27], inp_43d[27], nwaySelect_0n[43]);
  ND2 I2041 (nwayMuxOut_43n[28], inp_43d[28], nwaySelect_0n[43]);
  ND2 I2042 (nwayMuxOut_43n[29], inp_43d[29], nwaySelect_0n[43]);
  ND2 I2043 (nwayMuxOut_43n[30], inp_43d[30], nwaySelect_0n[43]);
  ND2 I2044 (nwayMuxOut_43n[31], inp_43d[31], nwaySelect_0n[43]);
  ND2 I2045 (nwayMuxOut_43n[32], inp_43d[32], nwaySelect_0n[43]);
  ND2 I2046 (nwayMuxOut_44n[0], inp_44d[0], nwaySelect_0n[44]);
  ND2 I2047 (nwayMuxOut_44n[1], inp_44d[1], nwaySelect_0n[44]);
  ND2 I2048 (nwayMuxOut_44n[2], inp_44d[2], nwaySelect_0n[44]);
  ND2 I2049 (nwayMuxOut_44n[3], inp_44d[3], nwaySelect_0n[44]);
  ND2 I2050 (nwayMuxOut_44n[4], inp_44d[4], nwaySelect_0n[44]);
  ND2 I2051 (nwayMuxOut_44n[5], inp_44d[5], nwaySelect_0n[44]);
  ND2 I2052 (nwayMuxOut_44n[6], inp_44d[6], nwaySelect_0n[44]);
  ND2 I2053 (nwayMuxOut_44n[7], inp_44d[7], nwaySelect_0n[44]);
  ND2 I2054 (nwayMuxOut_44n[8], inp_44d[8], nwaySelect_0n[44]);
  ND2 I2055 (nwayMuxOut_44n[9], inp_44d[9], nwaySelect_0n[44]);
  ND2 I2056 (nwayMuxOut_44n[10], inp_44d[10], nwaySelect_0n[44]);
  ND2 I2057 (nwayMuxOut_44n[11], inp_44d[11], nwaySelect_0n[44]);
  ND2 I2058 (nwayMuxOut_44n[12], inp_44d[12], nwaySelect_0n[44]);
  ND2 I2059 (nwayMuxOut_44n[13], inp_44d[13], nwaySelect_0n[44]);
  ND2 I2060 (nwayMuxOut_44n[14], inp_44d[14], nwaySelect_0n[44]);
  ND2 I2061 (nwayMuxOut_44n[15], inp_44d[15], nwaySelect_0n[44]);
  ND2 I2062 (nwayMuxOut_44n[16], inp_44d[16], nwaySelect_0n[44]);
  ND2 I2063 (nwayMuxOut_44n[17], inp_44d[17], nwaySelect_0n[44]);
  ND2 I2064 (nwayMuxOut_44n[18], inp_44d[18], nwaySelect_0n[44]);
  ND2 I2065 (nwayMuxOut_44n[19], inp_44d[19], nwaySelect_0n[44]);
  ND2 I2066 (nwayMuxOut_44n[20], inp_44d[20], nwaySelect_0n[44]);
  ND2 I2067 (nwayMuxOut_44n[21], inp_44d[21], nwaySelect_0n[44]);
  ND2 I2068 (nwayMuxOut_44n[22], inp_44d[22], nwaySelect_0n[44]);
  ND2 I2069 (nwayMuxOut_44n[23], inp_44d[23], nwaySelect_0n[44]);
  ND2 I2070 (nwayMuxOut_44n[24], inp_44d[24], nwaySelect_0n[44]);
  ND2 I2071 (nwayMuxOut_44n[25], inp_44d[25], nwaySelect_0n[44]);
  ND2 I2072 (nwayMuxOut_44n[26], inp_44d[26], nwaySelect_0n[44]);
  ND2 I2073 (nwayMuxOut_44n[27], inp_44d[27], nwaySelect_0n[44]);
  ND2 I2074 (nwayMuxOut_44n[28], inp_44d[28], nwaySelect_0n[44]);
  ND2 I2075 (nwayMuxOut_44n[29], inp_44d[29], nwaySelect_0n[44]);
  ND2 I2076 (nwayMuxOut_44n[30], inp_44d[30], nwaySelect_0n[44]);
  ND2 I2077 (nwayMuxOut_44n[31], inp_44d[31], nwaySelect_0n[44]);
  ND2 I2078 (nwayMuxOut_44n[32], inp_44d[32], nwaySelect_0n[44]);
  ND2 I2079 (nwayMuxOut_45n[0], inp_45d[0], nwaySelect_0n[45]);
  ND2 I2080 (nwayMuxOut_45n[1], inp_45d[1], nwaySelect_0n[45]);
  ND2 I2081 (nwayMuxOut_45n[2], inp_45d[2], nwaySelect_0n[45]);
  ND2 I2082 (nwayMuxOut_45n[3], inp_45d[3], nwaySelect_0n[45]);
  ND2 I2083 (nwayMuxOut_45n[4], inp_45d[4], nwaySelect_0n[45]);
  ND2 I2084 (nwayMuxOut_45n[5], inp_45d[5], nwaySelect_0n[45]);
  ND2 I2085 (nwayMuxOut_45n[6], inp_45d[6], nwaySelect_0n[45]);
  ND2 I2086 (nwayMuxOut_45n[7], inp_45d[7], nwaySelect_0n[45]);
  ND2 I2087 (nwayMuxOut_45n[8], inp_45d[8], nwaySelect_0n[45]);
  ND2 I2088 (nwayMuxOut_45n[9], inp_45d[9], nwaySelect_0n[45]);
  ND2 I2089 (nwayMuxOut_45n[10], inp_45d[10], nwaySelect_0n[45]);
  ND2 I2090 (nwayMuxOut_45n[11], inp_45d[11], nwaySelect_0n[45]);
  ND2 I2091 (nwayMuxOut_45n[12], inp_45d[12], nwaySelect_0n[45]);
  ND2 I2092 (nwayMuxOut_45n[13], inp_45d[13], nwaySelect_0n[45]);
  ND2 I2093 (nwayMuxOut_45n[14], inp_45d[14], nwaySelect_0n[45]);
  ND2 I2094 (nwayMuxOut_45n[15], inp_45d[15], nwaySelect_0n[45]);
  ND2 I2095 (nwayMuxOut_45n[16], inp_45d[16], nwaySelect_0n[45]);
  ND2 I2096 (nwayMuxOut_45n[17], inp_45d[17], nwaySelect_0n[45]);
  ND2 I2097 (nwayMuxOut_45n[18], inp_45d[18], nwaySelect_0n[45]);
  ND2 I2098 (nwayMuxOut_45n[19], inp_45d[19], nwaySelect_0n[45]);
  ND2 I2099 (nwayMuxOut_45n[20], inp_45d[20], nwaySelect_0n[45]);
  ND2 I2100 (nwayMuxOut_45n[21], inp_45d[21], nwaySelect_0n[45]);
  ND2 I2101 (nwayMuxOut_45n[22], inp_45d[22], nwaySelect_0n[45]);
  ND2 I2102 (nwayMuxOut_45n[23], inp_45d[23], nwaySelect_0n[45]);
  ND2 I2103 (nwayMuxOut_45n[24], inp_45d[24], nwaySelect_0n[45]);
  ND2 I2104 (nwayMuxOut_45n[25], inp_45d[25], nwaySelect_0n[45]);
  ND2 I2105 (nwayMuxOut_45n[26], inp_45d[26], nwaySelect_0n[45]);
  ND2 I2106 (nwayMuxOut_45n[27], inp_45d[27], nwaySelect_0n[45]);
  ND2 I2107 (nwayMuxOut_45n[28], inp_45d[28], nwaySelect_0n[45]);
  ND2 I2108 (nwayMuxOut_45n[29], inp_45d[29], nwaySelect_0n[45]);
  ND2 I2109 (nwayMuxOut_45n[30], inp_45d[30], nwaySelect_0n[45]);
  ND2 I2110 (nwayMuxOut_45n[31], inp_45d[31], nwaySelect_0n[45]);
  ND2 I2111 (nwayMuxOut_45n[32], inp_45d[32], nwaySelect_0n[45]);
  ND2 I2112 (nwayMuxOut_46n[0], inp_46d[0], nwaySelect_0n[46]);
  ND2 I2113 (nwayMuxOut_46n[1], inp_46d[1], nwaySelect_0n[46]);
  ND2 I2114 (nwayMuxOut_46n[2], inp_46d[2], nwaySelect_0n[46]);
  ND2 I2115 (nwayMuxOut_46n[3], inp_46d[3], nwaySelect_0n[46]);
  ND2 I2116 (nwayMuxOut_46n[4], inp_46d[4], nwaySelect_0n[46]);
  ND2 I2117 (nwayMuxOut_46n[5], inp_46d[5], nwaySelect_0n[46]);
  ND2 I2118 (nwayMuxOut_46n[6], inp_46d[6], nwaySelect_0n[46]);
  ND2 I2119 (nwayMuxOut_46n[7], inp_46d[7], nwaySelect_0n[46]);
  ND2 I2120 (nwayMuxOut_46n[8], inp_46d[8], nwaySelect_0n[46]);
  ND2 I2121 (nwayMuxOut_46n[9], inp_46d[9], nwaySelect_0n[46]);
  ND2 I2122 (nwayMuxOut_46n[10], inp_46d[10], nwaySelect_0n[46]);
  ND2 I2123 (nwayMuxOut_46n[11], inp_46d[11], nwaySelect_0n[46]);
  ND2 I2124 (nwayMuxOut_46n[12], inp_46d[12], nwaySelect_0n[46]);
  ND2 I2125 (nwayMuxOut_46n[13], inp_46d[13], nwaySelect_0n[46]);
  ND2 I2126 (nwayMuxOut_46n[14], inp_46d[14], nwaySelect_0n[46]);
  ND2 I2127 (nwayMuxOut_46n[15], inp_46d[15], nwaySelect_0n[46]);
  ND2 I2128 (nwayMuxOut_46n[16], inp_46d[16], nwaySelect_0n[46]);
  ND2 I2129 (nwayMuxOut_46n[17], inp_46d[17], nwaySelect_0n[46]);
  ND2 I2130 (nwayMuxOut_46n[18], inp_46d[18], nwaySelect_0n[46]);
  ND2 I2131 (nwayMuxOut_46n[19], inp_46d[19], nwaySelect_0n[46]);
  ND2 I2132 (nwayMuxOut_46n[20], inp_46d[20], nwaySelect_0n[46]);
  ND2 I2133 (nwayMuxOut_46n[21], inp_46d[21], nwaySelect_0n[46]);
  ND2 I2134 (nwayMuxOut_46n[22], inp_46d[22], nwaySelect_0n[46]);
  ND2 I2135 (nwayMuxOut_46n[23], inp_46d[23], nwaySelect_0n[46]);
  ND2 I2136 (nwayMuxOut_46n[24], inp_46d[24], nwaySelect_0n[46]);
  ND2 I2137 (nwayMuxOut_46n[25], inp_46d[25], nwaySelect_0n[46]);
  ND2 I2138 (nwayMuxOut_46n[26], inp_46d[26], nwaySelect_0n[46]);
  ND2 I2139 (nwayMuxOut_46n[27], inp_46d[27], nwaySelect_0n[46]);
  ND2 I2140 (nwayMuxOut_46n[28], inp_46d[28], nwaySelect_0n[46]);
  ND2 I2141 (nwayMuxOut_46n[29], inp_46d[29], nwaySelect_0n[46]);
  ND2 I2142 (nwayMuxOut_46n[30], inp_46d[30], nwaySelect_0n[46]);
  ND2 I2143 (nwayMuxOut_46n[31], inp_46d[31], nwaySelect_0n[46]);
  ND2 I2144 (nwayMuxOut_46n[32], inp_46d[32], nwaySelect_0n[46]);
  ND2 I2145 (nwayMuxOut_47n[0], inp_47d[0], nwaySelect_0n[47]);
  ND2 I2146 (nwayMuxOut_47n[1], inp_47d[1], nwaySelect_0n[47]);
  ND2 I2147 (nwayMuxOut_47n[2], inp_47d[2], nwaySelect_0n[47]);
  ND2 I2148 (nwayMuxOut_47n[3], inp_47d[3], nwaySelect_0n[47]);
  ND2 I2149 (nwayMuxOut_47n[4], inp_47d[4], nwaySelect_0n[47]);
  ND2 I2150 (nwayMuxOut_47n[5], inp_47d[5], nwaySelect_0n[47]);
  ND2 I2151 (nwayMuxOut_47n[6], inp_47d[6], nwaySelect_0n[47]);
  ND2 I2152 (nwayMuxOut_47n[7], inp_47d[7], nwaySelect_0n[47]);
  ND2 I2153 (nwayMuxOut_47n[8], inp_47d[8], nwaySelect_0n[47]);
  ND2 I2154 (nwayMuxOut_47n[9], inp_47d[9], nwaySelect_0n[47]);
  ND2 I2155 (nwayMuxOut_47n[10], inp_47d[10], nwaySelect_0n[47]);
  ND2 I2156 (nwayMuxOut_47n[11], inp_47d[11], nwaySelect_0n[47]);
  ND2 I2157 (nwayMuxOut_47n[12], inp_47d[12], nwaySelect_0n[47]);
  ND2 I2158 (nwayMuxOut_47n[13], inp_47d[13], nwaySelect_0n[47]);
  ND2 I2159 (nwayMuxOut_47n[14], inp_47d[14], nwaySelect_0n[47]);
  ND2 I2160 (nwayMuxOut_47n[15], inp_47d[15], nwaySelect_0n[47]);
  ND2 I2161 (nwayMuxOut_47n[16], inp_47d[16], nwaySelect_0n[47]);
  ND2 I2162 (nwayMuxOut_47n[17], inp_47d[17], nwaySelect_0n[47]);
  ND2 I2163 (nwayMuxOut_47n[18], inp_47d[18], nwaySelect_0n[47]);
  ND2 I2164 (nwayMuxOut_47n[19], inp_47d[19], nwaySelect_0n[47]);
  ND2 I2165 (nwayMuxOut_47n[20], inp_47d[20], nwaySelect_0n[47]);
  ND2 I2166 (nwayMuxOut_47n[21], inp_47d[21], nwaySelect_0n[47]);
  ND2 I2167 (nwayMuxOut_47n[22], inp_47d[22], nwaySelect_0n[47]);
  ND2 I2168 (nwayMuxOut_47n[23], inp_47d[23], nwaySelect_0n[47]);
  ND2 I2169 (nwayMuxOut_47n[24], inp_47d[24], nwaySelect_0n[47]);
  ND2 I2170 (nwayMuxOut_47n[25], inp_47d[25], nwaySelect_0n[47]);
  ND2 I2171 (nwayMuxOut_47n[26], inp_47d[26], nwaySelect_0n[47]);
  ND2 I2172 (nwayMuxOut_47n[27], inp_47d[27], nwaySelect_0n[47]);
  ND2 I2173 (nwayMuxOut_47n[28], inp_47d[28], nwaySelect_0n[47]);
  ND2 I2174 (nwayMuxOut_47n[29], inp_47d[29], nwaySelect_0n[47]);
  ND2 I2175 (nwayMuxOut_47n[30], inp_47d[30], nwaySelect_0n[47]);
  ND2 I2176 (nwayMuxOut_47n[31], inp_47d[31], nwaySelect_0n[47]);
  ND2 I2177 (nwayMuxOut_47n[32], inp_47d[32], nwaySelect_0n[47]);
  ND2 I2178 (nwayMuxOut_48n[0], inp_48d[0], nwaySelect_0n[48]);
  ND2 I2179 (nwayMuxOut_48n[1], inp_48d[1], nwaySelect_0n[48]);
  ND2 I2180 (nwayMuxOut_48n[2], inp_48d[2], nwaySelect_0n[48]);
  ND2 I2181 (nwayMuxOut_48n[3], inp_48d[3], nwaySelect_0n[48]);
  ND2 I2182 (nwayMuxOut_48n[4], inp_48d[4], nwaySelect_0n[48]);
  ND2 I2183 (nwayMuxOut_48n[5], inp_48d[5], nwaySelect_0n[48]);
  ND2 I2184 (nwayMuxOut_48n[6], inp_48d[6], nwaySelect_0n[48]);
  ND2 I2185 (nwayMuxOut_48n[7], inp_48d[7], nwaySelect_0n[48]);
  ND2 I2186 (nwayMuxOut_48n[8], inp_48d[8], nwaySelect_0n[48]);
  ND2 I2187 (nwayMuxOut_48n[9], inp_48d[9], nwaySelect_0n[48]);
  ND2 I2188 (nwayMuxOut_48n[10], inp_48d[10], nwaySelect_0n[48]);
  ND2 I2189 (nwayMuxOut_48n[11], inp_48d[11], nwaySelect_0n[48]);
  ND2 I2190 (nwayMuxOut_48n[12], inp_48d[12], nwaySelect_0n[48]);
  ND2 I2191 (nwayMuxOut_48n[13], inp_48d[13], nwaySelect_0n[48]);
  ND2 I2192 (nwayMuxOut_48n[14], inp_48d[14], nwaySelect_0n[48]);
  ND2 I2193 (nwayMuxOut_48n[15], inp_48d[15], nwaySelect_0n[48]);
  ND2 I2194 (nwayMuxOut_48n[16], inp_48d[16], nwaySelect_0n[48]);
  ND2 I2195 (nwayMuxOut_48n[17], inp_48d[17], nwaySelect_0n[48]);
  ND2 I2196 (nwayMuxOut_48n[18], inp_48d[18], nwaySelect_0n[48]);
  ND2 I2197 (nwayMuxOut_48n[19], inp_48d[19], nwaySelect_0n[48]);
  ND2 I2198 (nwayMuxOut_48n[20], inp_48d[20], nwaySelect_0n[48]);
  ND2 I2199 (nwayMuxOut_48n[21], inp_48d[21], nwaySelect_0n[48]);
  ND2 I2200 (nwayMuxOut_48n[22], inp_48d[22], nwaySelect_0n[48]);
  ND2 I2201 (nwayMuxOut_48n[23], inp_48d[23], nwaySelect_0n[48]);
  ND2 I2202 (nwayMuxOut_48n[24], inp_48d[24], nwaySelect_0n[48]);
  ND2 I2203 (nwayMuxOut_48n[25], inp_48d[25], nwaySelect_0n[48]);
  ND2 I2204 (nwayMuxOut_48n[26], inp_48d[26], nwaySelect_0n[48]);
  ND2 I2205 (nwayMuxOut_48n[27], inp_48d[27], nwaySelect_0n[48]);
  ND2 I2206 (nwayMuxOut_48n[28], inp_48d[28], nwaySelect_0n[48]);
  ND2 I2207 (nwayMuxOut_48n[29], inp_48d[29], nwaySelect_0n[48]);
  ND2 I2208 (nwayMuxOut_48n[30], inp_48d[30], nwaySelect_0n[48]);
  ND2 I2209 (nwayMuxOut_48n[31], inp_48d[31], nwaySelect_0n[48]);
  ND2 I2210 (nwayMuxOut_48n[32], inp_48d[32], nwaySelect_0n[48]);
  OR2 I2211 (nwaySelect_0n[0], inp_0a, inp_0r);
  OR2 I2212 (nwaySelect_0n[1], inp_1a, inp_1r);
  OR2 I2213 (nwaySelect_0n[2], inp_2a, inp_2r);
  OR2 I2214 (nwaySelect_0n[3], inp_3a, inp_3r);
  OR2 I2215 (nwaySelect_0n[4], inp_4a, inp_4r);
  OR2 I2216 (nwaySelect_0n[5], inp_5a, inp_5r);
  OR2 I2217 (nwaySelect_0n[6], inp_6a, inp_6r);
  OR2 I2218 (nwaySelect_0n[7], inp_7a, inp_7r);
  OR2 I2219 (nwaySelect_0n[8], inp_8a, inp_8r);
  OR2 I2220 (nwaySelect_0n[9], inp_9a, inp_9r);
  OR2 I2221 (nwaySelect_0n[10], inp_10a, inp_10r);
  OR2 I2222 (nwaySelect_0n[11], inp_11a, inp_11r);
  OR2 I2223 (nwaySelect_0n[12], inp_12a, inp_12r);
  OR2 I2224 (nwaySelect_0n[13], inp_13a, inp_13r);
  OR2 I2225 (nwaySelect_0n[14], inp_14a, inp_14r);
  OR2 I2226 (nwaySelect_0n[15], inp_15a, inp_15r);
  OR2 I2227 (nwaySelect_0n[16], inp_16a, inp_16r);
  OR2 I2228 (nwaySelect_0n[17], inp_17a, inp_17r);
  OR2 I2229 (nwaySelect_0n[18], inp_18a, inp_18r);
  OR2 I2230 (nwaySelect_0n[19], inp_19a, inp_19r);
  OR2 I2231 (nwaySelect_0n[20], inp_20a, inp_20r);
  OR2 I2232 (nwaySelect_0n[21], inp_21a, inp_21r);
  OR2 I2233 (nwaySelect_0n[22], inp_22a, inp_22r);
  OR2 I2234 (nwaySelect_0n[23], inp_23a, inp_23r);
  OR2 I2235 (nwaySelect_0n[24], inp_24a, inp_24r);
  OR2 I2236 (nwaySelect_0n[25], inp_25a, inp_25r);
  OR2 I2237 (nwaySelect_0n[26], inp_26a, inp_26r);
  OR2 I2238 (nwaySelect_0n[27], inp_27a, inp_27r);
  OR2 I2239 (nwaySelect_0n[28], inp_28a, inp_28r);
  OR2 I2240 (nwaySelect_0n[29], inp_29a, inp_29r);
  OR2 I2241 (nwaySelect_0n[30], inp_30a, inp_30r);
  OR2 I2242 (nwaySelect_0n[31], inp_31a, inp_31r);
  OR2 I2243 (nwaySelect_0n[32], inp_32a, inp_32r);
  OR2 I2244 (nwaySelect_0n[33], inp_33a, inp_33r);
  OR2 I2245 (nwaySelect_0n[34], inp_34a, inp_34r);
  OR2 I2246 (nwaySelect_0n[35], inp_35a, inp_35r);
  OR2 I2247 (nwaySelect_0n[36], inp_36a, inp_36r);
  OR2 I2248 (nwaySelect_0n[37], inp_37a, inp_37r);
  OR2 I2249 (nwaySelect_0n[38], inp_38a, inp_38r);
  OR2 I2250 (nwaySelect_0n[39], inp_39a, inp_39r);
  OR2 I2251 (nwaySelect_0n[40], inp_40a, inp_40r);
  OR2 I2252 (nwaySelect_0n[41], inp_41a, inp_41r);
  OR2 I2253 (nwaySelect_0n[42], inp_42a, inp_42r);
  OR2 I2254 (nwaySelect_0n[43], inp_43a, inp_43r);
  OR2 I2255 (nwaySelect_0n[44], inp_44a, inp_44r);
  OR2 I2256 (nwaySelect_0n[45], inp_45a, inp_45r);
  OR2 I2257 (nwaySelect_0n[46], inp_46a, inp_46r);
  OR2 I2258 (nwaySelect_0n[47], inp_47a, inp_47r);
  OR2 I2259 (nwaySelect_0n[48], inp_48a, inp_48r);
  C2 I2260 (inp_0a, inp_0r, out_0a);
  C2 I2261 (inp_1a, inp_1r, out_0a);
  C2 I2262 (inp_2a, inp_2r, out_0a);
  C2 I2263 (inp_3a, inp_3r, out_0a);
  C2 I2264 (inp_4a, inp_4r, out_0a);
  C2 I2265 (inp_5a, inp_5r, out_0a);
  C2 I2266 (inp_6a, inp_6r, out_0a);
  C2 I2267 (inp_7a, inp_7r, out_0a);
  C2 I2268 (inp_8a, inp_8r, out_0a);
  C2 I2269 (inp_9a, inp_9r, out_0a);
  C2 I2270 (inp_10a, inp_10r, out_0a);
  C2 I2271 (inp_11a, inp_11r, out_0a);
  C2 I2272 (inp_12a, inp_12r, out_0a);
  C2 I2273 (inp_13a, inp_13r, out_0a);
  C2 I2274 (inp_14a, inp_14r, out_0a);
  C2 I2275 (inp_15a, inp_15r, out_0a);
  C2 I2276 (inp_16a, inp_16r, out_0a);
  C2 I2277 (inp_17a, inp_17r, out_0a);
  C2 I2278 (inp_18a, inp_18r, out_0a);
  C2 I2279 (inp_19a, inp_19r, out_0a);
  C2 I2280 (inp_20a, inp_20r, out_0a);
  C2 I2281 (inp_21a, inp_21r, out_0a);
  C2 I2282 (inp_22a, inp_22r, out_0a);
  C2 I2283 (inp_23a, inp_23r, out_0a);
  C2 I2284 (inp_24a, inp_24r, out_0a);
  C2 I2285 (inp_25a, inp_25r, out_0a);
  C2 I2286 (inp_26a, inp_26r, out_0a);
  C2 I2287 (inp_27a, inp_27r, out_0a);
  C2 I2288 (inp_28a, inp_28r, out_0a);
  C2 I2289 (inp_29a, inp_29r, out_0a);
  C2 I2290 (inp_30a, inp_30r, out_0a);
  C2 I2291 (inp_31a, inp_31r, out_0a);
  C2 I2292 (inp_32a, inp_32r, out_0a);
  C2 I2293 (inp_33a, inp_33r, out_0a);
  C2 I2294 (inp_34a, inp_34r, out_0a);
  C2 I2295 (inp_35a, inp_35r, out_0a);
  C2 I2296 (inp_36a, inp_36r, out_0a);
  C2 I2297 (inp_37a, inp_37r, out_0a);
  C2 I2298 (inp_38a, inp_38r, out_0a);
  C2 I2299 (inp_39a, inp_39r, out_0a);
  C2 I2300 (inp_40a, inp_40r, out_0a);
  C2 I2301 (inp_41a, inp_41r, out_0a);
  C2 I2302 (inp_42a, inp_42r, out_0a);
  C2 I2303 (inp_43a, inp_43r, out_0a);
  C2 I2304 (inp_44a, inp_44r, out_0a);
  C2 I2305 (inp_45a, inp_45r, out_0a);
  C2 I2306 (inp_46a, inp_46r, out_0a);
  C2 I2307 (inp_47a, inp_47r, out_0a);
  C2 I2308 (inp_48a, inp_48r, out_0a);
  NR4 I2309 (internal_0n[561], inp_0r, inp_1r, inp_2r, inp_3r);
  NR4 I2310 (internal_0n[562], inp_4r, inp_5r, inp_6r, inp_7r);
  NR4 I2311 (internal_0n[563], inp_8r, inp_9r, inp_10r, inp_11r);
  NR4 I2312 (internal_0n[564], inp_12r, inp_13r, inp_14r, inp_15r);
  NR4 I2313 (internal_0n[565], inp_16r, inp_17r, inp_18r, inp_19r);
  NR4 I2314 (internal_0n[566], inp_20r, inp_21r, inp_22r, inp_23r);
  NR4 I2315 (internal_0n[567], inp_24r, inp_25r, inp_26r, inp_27r);
  NR4 I2316 (internal_0n[568], inp_28r, inp_29r, inp_30r, inp_31r);
  NR4 I2317 (internal_0n[569], inp_32r, inp_33r, inp_34r, inp_35r);
  NR4 I2318 (internal_0n[570], inp_36r, inp_37r, inp_38r, inp_39r);
  NR4 I2319 (internal_0n[571], inp_40r, inp_41r, inp_42r, inp_43r);
  NR2 I2320 (internal_0n[572], inp_44r, inp_45r);
  NR3 I2321 (internal_0n[573], inp_46r, inp_47r, inp_48r);
  ND4 I2322 (internal_0n[574], internal_0n[561], internal_0n[562], internal_0n[563], internal_0n[564]);
  ND4 I2323 (internal_0n[575], internal_0n[565], internal_0n[566], internal_0n[567], internal_0n[568]);
  ND2 I2324 (internal_0n[576], internal_0n[569], internal_0n[570]);
  ND3 I2325 (internal_0n[577], internal_0n[571], internal_0n[572], internal_0n[573]);
  OR4 I2326 (out_0r, internal_0n[574], internal_0n[575], internal_0n[576], internal_0n[577]);
endmodule

module BrzCase_1_2_s5_0_3b1 (
  inp_0r, inp_0a, inp_0d,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a
);
  input inp_0r;
  output inp_0a;
  input inp_0d;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  wire t_0n;
  wire c_0n;
  wire elseAck_0n;
  wire [1:0] int0_0n;
  OR2 I0 (inp_0a, activateOut_0a, activateOut_1a);
  assign int0_0n[0] = c_0n;
  assign int0_0n[1] = t_0n;
  assign activateOut_1r = int0_0n[1];
  assign activateOut_0r = int0_0n[0];
  demux2 I5 (inp_0r, c_0n, t_0n, inp_0d);
endmodule

module BrzCombine_17_1_16 (
  out_0r, out_0a, out_0d,
  LSInp_0r, LSInp_0a, LSInp_0d,
  MSInp_0r, MSInp_0a, MSInp_0d
);
  input out_0r;
  output out_0a;
  output [16:0] out_0d;
  output LSInp_0r;
  input LSInp_0a;
  input LSInp_0d;
  output MSInp_0r;
  input MSInp_0a;
  input [15:0] MSInp_0d;
  C2 I0 (out_0a, LSInp_0a, MSInp_0a);
  assign LSInp_0r = out_0r;
  assign MSInp_0r = out_0r;
  assign out_0d[0] = LSInp_0d;
  assign out_0d[1] = MSInp_0d[0];
  assign out_0d[2] = MSInp_0d[1];
  assign out_0d[3] = MSInp_0d[2];
  assign out_0d[4] = MSInp_0d[3];
  assign out_0d[5] = MSInp_0d[4];
  assign out_0d[6] = MSInp_0d[5];
  assign out_0d[7] = MSInp_0d[6];
  assign out_0d[8] = MSInp_0d[7];
  assign out_0d[9] = MSInp_0d[8];
  assign out_0d[10] = MSInp_0d[9];
  assign out_0d[11] = MSInp_0d[10];
  assign out_0d[12] = MSInp_0d[11];
  assign out_0d[13] = MSInp_0d[12];
  assign out_0d[14] = MSInp_0d[13];
  assign out_0d[15] = MSInp_0d[14];
  assign out_0d[16] = MSInp_0d[15];
endmodule

module BrzCombine_33_17_16 (
  out_0r, out_0a, out_0d,
  LSInp_0r, LSInp_0a, LSInp_0d,
  MSInp_0r, MSInp_0a, MSInp_0d
);
  input out_0r;
  output out_0a;
  output [32:0] out_0d;
  output LSInp_0r;
  input LSInp_0a;
  input [16:0] LSInp_0d;
  output MSInp_0r;
  input MSInp_0a;
  input [15:0] MSInp_0d;
  C2 I0 (out_0a, LSInp_0a, MSInp_0a);
  assign LSInp_0r = out_0r;
  assign MSInp_0r = out_0r;
  assign out_0d[0] = LSInp_0d[0];
  assign out_0d[1] = LSInp_0d[1];
  assign out_0d[2] = LSInp_0d[2];
  assign out_0d[3] = LSInp_0d[3];
  assign out_0d[4] = LSInp_0d[4];
  assign out_0d[5] = LSInp_0d[5];
  assign out_0d[6] = LSInp_0d[6];
  assign out_0d[7] = LSInp_0d[7];
  assign out_0d[8] = LSInp_0d[8];
  assign out_0d[9] = LSInp_0d[9];
  assign out_0d[10] = LSInp_0d[10];
  assign out_0d[11] = LSInp_0d[11];
  assign out_0d[12] = LSInp_0d[12];
  assign out_0d[13] = LSInp_0d[13];
  assign out_0d[14] = LSInp_0d[14];
  assign out_0d[15] = LSInp_0d[15];
  assign out_0d[16] = LSInp_0d[16];
  assign out_0d[17] = MSInp_0d[0];
  assign out_0d[18] = MSInp_0d[1];
  assign out_0d[19] = MSInp_0d[2];
  assign out_0d[20] = MSInp_0d[3];
  assign out_0d[21] = MSInp_0d[4];
  assign out_0d[22] = MSInp_0d[5];
  assign out_0d[23] = MSInp_0d[6];
  assign out_0d[24] = MSInp_0d[7];
  assign out_0d[25] = MSInp_0d[8];
  assign out_0d[26] = MSInp_0d[9];
  assign out_0d[27] = MSInp_0d[10];
  assign out_0d[28] = MSInp_0d[11];
  assign out_0d[29] = MSInp_0d[12];
  assign out_0d[30] = MSInp_0d[13];
  assign out_0d[31] = MSInp_0d[14];
  assign out_0d[32] = MSInp_0d[15];
endmodule

module BrzCombine_33_32_1 (
  out_0r, out_0a, out_0d,
  LSInp_0r, LSInp_0a, LSInp_0d,
  MSInp_0r, MSInp_0a, MSInp_0d
);
  input out_0r;
  output out_0a;
  output [32:0] out_0d;
  output LSInp_0r;
  input LSInp_0a;
  input [31:0] LSInp_0d;
  output MSInp_0r;
  input MSInp_0a;
  input MSInp_0d;
  C2 I0 (out_0a, LSInp_0a, MSInp_0a);
  assign LSInp_0r = out_0r;
  assign MSInp_0r = out_0r;
  assign out_0d[0] = LSInp_0d[0];
  assign out_0d[1] = LSInp_0d[1];
  assign out_0d[2] = LSInp_0d[2];
  assign out_0d[3] = LSInp_0d[3];
  assign out_0d[4] = LSInp_0d[4];
  assign out_0d[5] = LSInp_0d[5];
  assign out_0d[6] = LSInp_0d[6];
  assign out_0d[7] = LSInp_0d[7];
  assign out_0d[8] = LSInp_0d[8];
  assign out_0d[9] = LSInp_0d[9];
  assign out_0d[10] = LSInp_0d[10];
  assign out_0d[11] = LSInp_0d[11];
  assign out_0d[12] = LSInp_0d[12];
  assign out_0d[13] = LSInp_0d[13];
  assign out_0d[14] = LSInp_0d[14];
  assign out_0d[15] = LSInp_0d[15];
  assign out_0d[16] = LSInp_0d[16];
  assign out_0d[17] = LSInp_0d[17];
  assign out_0d[18] = LSInp_0d[18];
  assign out_0d[19] = LSInp_0d[19];
  assign out_0d[20] = LSInp_0d[20];
  assign out_0d[21] = LSInp_0d[21];
  assign out_0d[22] = LSInp_0d[22];
  assign out_0d[23] = LSInp_0d[23];
  assign out_0d[24] = LSInp_0d[24];
  assign out_0d[25] = LSInp_0d[25];
  assign out_0d[26] = LSInp_0d[26];
  assign out_0d[27] = LSInp_0d[27];
  assign out_0d[28] = LSInp_0d[28];
  assign out_0d[29] = LSInp_0d[29];
  assign out_0d[30] = LSInp_0d[30];
  assign out_0d[31] = LSInp_0d[31];
  assign out_0d[32] = MSInp_0d;
endmodule

module telem (
  Ar,
  Aa,
  Br,
  Ba
);
  input Ar;
  output Aa;
  output Br;
  input Ba;
  wire s_0n;
  ACU0D1 I0 (Aa, Ba, Ar);
  IV I1 (s_0n, Aa);
  AN2 I2 (Br, Ar, s_0n);
endmodule

module BrzConcur_2 (
  activate_0r, activate_0a,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a
);
  input activate_0r;
  output activate_0a;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  wire [1:0] acks_0n;
  C2 I0 (activate_0a, acks_0n[0], acks_0n[1]);
  telem I1 (activate_0r, acks_0n[0], activateOut_0r, activateOut_0a);
  telem I2 (activate_0r, acks_0n[1], activateOut_1r, activateOut_1a);
endmodule

module BrzConcur_3 (
  activate_0r, activate_0a,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a,
  activateOut_2r, activateOut_2a
);
  input activate_0r;
  output activate_0a;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  output activateOut_2r;
  input activateOut_2a;
  wire [2:0] acks_0n;
  C3 I0 (activate_0a, acks_0n[0], acks_0n[1], acks_0n[2]);
  telem I1 (activate_0r, acks_0n[0], activateOut_0r, activateOut_0a);
  telem I2 (activate_0r, acks_0n[1], activateOut_1r, activateOut_1a);
  telem I3 (activate_0r, acks_0n[2], activateOut_2r, activateOut_2a);
endmodule

module BrzConstant_1_0 (
  out_0r, out_0a, out_0d
);
  input out_0r;
  output out_0a;
  output out_0d;
  wire gnd;
  GND gnd_cell_instance (gnd);
  assign out_0a = out_0r;
  assign out_0d = gnd;
endmodule

module BrzConstant_17_0 (
  out_0r, out_0a, out_0d
);
  input out_0r;
  output out_0a;
  output [16:0] out_0d;
  wire gnd;
  GND gnd_cell_instance (gnd);
  assign out_0a = out_0r;
  assign out_0d[0] = gnd;
  assign out_0d[1] = gnd;
  assign out_0d[2] = gnd;
  assign out_0d[3] = gnd;
  assign out_0d[4] = gnd;
  assign out_0d[5] = gnd;
  assign out_0d[6] = gnd;
  assign out_0d[7] = gnd;
  assign out_0d[8] = gnd;
  assign out_0d[9] = gnd;
  assign out_0d[10] = gnd;
  assign out_0d[11] = gnd;
  assign out_0d[12] = gnd;
  assign out_0d[13] = gnd;
  assign out_0d[14] = gnd;
  assign out_0d[15] = gnd;
  assign out_0d[16] = gnd;
endmodule

module BrzFetch_1_s5_false (
  activate_0r, activate_0a,
  inp_0r, inp_0a, inp_0d,
  out_0r, out_0a, out_0d
);
  input activate_0r;
  output activate_0a;
  output inp_0r;
  input inp_0a;
  input inp_0d;
  output out_0r;
  input out_0a;
  output out_0d;
  assign activate_0a = out_0a;
  assign out_0r = inp_0a;
  assign inp_0r = activate_0r;
  assign out_0d = inp_0d;
endmodule

module BrzFetch_16_s5_false (
  activate_0r, activate_0a,
  inp_0r, inp_0a, inp_0d,
  out_0r, out_0a, out_0d
);
  input activate_0r;
  output activate_0a;
  output inp_0r;
  input inp_0a;
  input [15:0] inp_0d;
  output out_0r;
  input out_0a;
  output [15:0] out_0d;
  assign activate_0a = out_0a;
  assign out_0r = inp_0a;
  assign inp_0r = activate_0r;
  assign out_0d[0] = inp_0d[0];
  assign out_0d[1] = inp_0d[1];
  assign out_0d[2] = inp_0d[2];
  assign out_0d[3] = inp_0d[3];
  assign out_0d[4] = inp_0d[4];
  assign out_0d[5] = inp_0d[5];
  assign out_0d[6] = inp_0d[6];
  assign out_0d[7] = inp_0d[7];
  assign out_0d[8] = inp_0d[8];
  assign out_0d[9] = inp_0d[9];
  assign out_0d[10] = inp_0d[10];
  assign out_0d[11] = inp_0d[11];
  assign out_0d[12] = inp_0d[12];
  assign out_0d[13] = inp_0d[13];
  assign out_0d[14] = inp_0d[14];
  assign out_0d[15] = inp_0d[15];
endmodule

module BrzFetch_32_s5_false (
  activate_0r, activate_0a,
  inp_0r, inp_0a, inp_0d,
  out_0r, out_0a, out_0d
);
  input activate_0r;
  output activate_0a;
  output inp_0r;
  input inp_0a;
  input [31:0] inp_0d;
  output out_0r;
  input out_0a;
  output [31:0] out_0d;
  assign activate_0a = out_0a;
  assign out_0r = inp_0a;
  assign inp_0r = activate_0r;
  assign out_0d[0] = inp_0d[0];
  assign out_0d[1] = inp_0d[1];
  assign out_0d[2] = inp_0d[2];
  assign out_0d[3] = inp_0d[3];
  assign out_0d[4] = inp_0d[4];
  assign out_0d[5] = inp_0d[5];
  assign out_0d[6] = inp_0d[6];
  assign out_0d[7] = inp_0d[7];
  assign out_0d[8] = inp_0d[8];
  assign out_0d[9] = inp_0d[9];
  assign out_0d[10] = inp_0d[10];
  assign out_0d[11] = inp_0d[11];
  assign out_0d[12] = inp_0d[12];
  assign out_0d[13] = inp_0d[13];
  assign out_0d[14] = inp_0d[14];
  assign out_0d[15] = inp_0d[15];
  assign out_0d[16] = inp_0d[16];
  assign out_0d[17] = inp_0d[17];
  assign out_0d[18] = inp_0d[18];
  assign out_0d[19] = inp_0d[19];
  assign out_0d[20] = inp_0d[20];
  assign out_0d[21] = inp_0d[21];
  assign out_0d[22] = inp_0d[22];
  assign out_0d[23] = inp_0d[23];
  assign out_0d[24] = inp_0d[24];
  assign out_0d[25] = inp_0d[25];
  assign out_0d[26] = inp_0d[26];
  assign out_0d[27] = inp_0d[27];
  assign out_0d[28] = inp_0d[28];
  assign out_0d[29] = inp_0d[29];
  assign out_0d[30] = inp_0d[30];
  assign out_0d[31] = inp_0d[31];
endmodule

module BrzFetch_33_s5_false (
  activate_0r, activate_0a,
  inp_0r, inp_0a, inp_0d,
  out_0r, out_0a, out_0d
);
  input activate_0r;
  output activate_0a;
  output inp_0r;
  input inp_0a;
  input [32:0] inp_0d;
  output out_0r;
  input out_0a;
  output [32:0] out_0d;
  assign activate_0a = out_0a;
  assign out_0r = inp_0a;
  assign inp_0r = activate_0r;
  assign out_0d[0] = inp_0d[0];
  assign out_0d[1] = inp_0d[1];
  assign out_0d[2] = inp_0d[2];
  assign out_0d[3] = inp_0d[3];
  assign out_0d[4] = inp_0d[4];
  assign out_0d[5] = inp_0d[5];
  assign out_0d[6] = inp_0d[6];
  assign out_0d[7] = inp_0d[7];
  assign out_0d[8] = inp_0d[8];
  assign out_0d[9] = inp_0d[9];
  assign out_0d[10] = inp_0d[10];
  assign out_0d[11] = inp_0d[11];
  assign out_0d[12] = inp_0d[12];
  assign out_0d[13] = inp_0d[13];
  assign out_0d[14] = inp_0d[14];
  assign out_0d[15] = inp_0d[15];
  assign out_0d[16] = inp_0d[16];
  assign out_0d[17] = inp_0d[17];
  assign out_0d[18] = inp_0d[18];
  assign out_0d[19] = inp_0d[19];
  assign out_0d[20] = inp_0d[20];
  assign out_0d[21] = inp_0d[21];
  assign out_0d[22] = inp_0d[22];
  assign out_0d[23] = inp_0d[23];
  assign out_0d[24] = inp_0d[24];
  assign out_0d[25] = inp_0d[25];
  assign out_0d[26] = inp_0d[26];
  assign out_0d[27] = inp_0d[27];
  assign out_0d[28] = inp_0d[28];
  assign out_0d[29] = inp_0d[29];
  assign out_0d[30] = inp_0d[30];
  assign out_0d[31] = inp_0d[31];
  assign out_0d[32] = inp_0d[32];
endmodule

module BrzLoop (
  activate_0r, activate_0a,
  activateOut_0r, activateOut_0a
);
  input activate_0r;
  output activate_0a;
  output activateOut_0r;
  input activateOut_0a;
  wire nReq_0n;
  wire gnd;
  GND gnd_cell_instance (gnd);
  IV I0 (nReq_0n, activate_0r);
  NR2 I1 (activateOut_0r, nReq_0n, activateOut_0a);
  assign activate_0a = gnd;
endmodule

module selem (
  Ar,
  Aa,
  Br,
  Ba
);
  input Ar;
  output Aa;
  output Br;
  input Ba;
  wire s_0n;
  NC2P I0 (s_0n, Ar, Ba);
  NR2 I1 (Aa, Ba, s_0n);
  AN2 I2 (Br, Ar, s_0n);
endmodule

module BrzSequence_2_s1_S (
  activate_0r, activate_0a,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a
);
  input activate_0r;
  output activate_0a;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  wire [1:0] sreq_0n;
  assign activate_0a = activateOut_1a;
  assign activateOut_1r = sreq_0n[1];
  assign sreq_0n[0] = activate_0r;
  selem I3 (sreq_0n[0], sreq_0n[1], activateOut_0r, activateOut_0a);
endmodule

module BrzSequence_35_s34_SSSSSSSSSSSSSSSSSSSSSSS_m3m (
  activate_0r, activate_0a,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a,
  activateOut_2r, activateOut_2a,
  activateOut_3r, activateOut_3a,
  activateOut_4r, activateOut_4a,
  activateOut_5r, activateOut_5a,
  activateOut_6r, activateOut_6a,
  activateOut_7r, activateOut_7a,
  activateOut_8r, activateOut_8a,
  activateOut_9r, activateOut_9a,
  activateOut_10r, activateOut_10a,
  activateOut_11r, activateOut_11a,
  activateOut_12r, activateOut_12a,
  activateOut_13r, activateOut_13a,
  activateOut_14r, activateOut_14a,
  activateOut_15r, activateOut_15a,
  activateOut_16r, activateOut_16a,
  activateOut_17r, activateOut_17a,
  activateOut_18r, activateOut_18a,
  activateOut_19r, activateOut_19a,
  activateOut_20r, activateOut_20a,
  activateOut_21r, activateOut_21a,
  activateOut_22r, activateOut_22a,
  activateOut_23r, activateOut_23a,
  activateOut_24r, activateOut_24a,
  activateOut_25r, activateOut_25a,
  activateOut_26r, activateOut_26a,
  activateOut_27r, activateOut_27a,
  activateOut_28r, activateOut_28a,
  activateOut_29r, activateOut_29a,
  activateOut_30r, activateOut_30a,
  activateOut_31r, activateOut_31a,
  activateOut_32r, activateOut_32a,
  activateOut_33r, activateOut_33a,
  activateOut_34r, activateOut_34a
);
  input activate_0r;
  output activate_0a;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  output activateOut_2r;
  input activateOut_2a;
  output activateOut_3r;
  input activateOut_3a;
  output activateOut_4r;
  input activateOut_4a;
  output activateOut_5r;
  input activateOut_5a;
  output activateOut_6r;
  input activateOut_6a;
  output activateOut_7r;
  input activateOut_7a;
  output activateOut_8r;
  input activateOut_8a;
  output activateOut_9r;
  input activateOut_9a;
  output activateOut_10r;
  input activateOut_10a;
  output activateOut_11r;
  input activateOut_11a;
  output activateOut_12r;
  input activateOut_12a;
  output activateOut_13r;
  input activateOut_13a;
  output activateOut_14r;
  input activateOut_14a;
  output activateOut_15r;
  input activateOut_15a;
  output activateOut_16r;
  input activateOut_16a;
  output activateOut_17r;
  input activateOut_17a;
  output activateOut_18r;
  input activateOut_18a;
  output activateOut_19r;
  input activateOut_19a;
  output activateOut_20r;
  input activateOut_20a;
  output activateOut_21r;
  input activateOut_21a;
  output activateOut_22r;
  input activateOut_22a;
  output activateOut_23r;
  input activateOut_23a;
  output activateOut_24r;
  input activateOut_24a;
  output activateOut_25r;
  input activateOut_25a;
  output activateOut_26r;
  input activateOut_26a;
  output activateOut_27r;
  input activateOut_27a;
  output activateOut_28r;
  input activateOut_28a;
  output activateOut_29r;
  input activateOut_29a;
  output activateOut_30r;
  input activateOut_30a;
  output activateOut_31r;
  input activateOut_31a;
  output activateOut_32r;
  input activateOut_32a;
  output activateOut_33r;
  input activateOut_33a;
  output activateOut_34r;
  input activateOut_34a;
  wire [34:0] sreq_0n;
  assign activate_0a = activateOut_34a;
  assign activateOut_34r = sreq_0n[34];
  assign sreq_0n[0] = activate_0r;
  selem I3 (sreq_0n[33], sreq_0n[34], activateOut_33r, activateOut_33a);
  selem I4 (sreq_0n[32], sreq_0n[33], activateOut_32r, activateOut_32a);
  selem I5 (sreq_0n[31], sreq_0n[32], activateOut_31r, activateOut_31a);
  selem I6 (sreq_0n[30], sreq_0n[31], activateOut_30r, activateOut_30a);
  selem I7 (sreq_0n[29], sreq_0n[30], activateOut_29r, activateOut_29a);
  selem I8 (sreq_0n[28], sreq_0n[29], activateOut_28r, activateOut_28a);
  selem I9 (sreq_0n[27], sreq_0n[28], activateOut_27r, activateOut_27a);
  selem I10 (sreq_0n[26], sreq_0n[27], activateOut_26r, activateOut_26a);
  selem I11 (sreq_0n[25], sreq_0n[26], activateOut_25r, activateOut_25a);
  selem I12 (sreq_0n[24], sreq_0n[25], activateOut_24r, activateOut_24a);
  selem I13 (sreq_0n[23], sreq_0n[24], activateOut_23r, activateOut_23a);
  selem I14 (sreq_0n[22], sreq_0n[23], activateOut_22r, activateOut_22a);
  selem I15 (sreq_0n[21], sreq_0n[22], activateOut_21r, activateOut_21a);
  selem I16 (sreq_0n[20], sreq_0n[21], activateOut_20r, activateOut_20a);
  selem I17 (sreq_0n[19], sreq_0n[20], activateOut_19r, activateOut_19a);
  selem I18 (sreq_0n[18], sreq_0n[19], activateOut_18r, activateOut_18a);
  selem I19 (sreq_0n[17], sreq_0n[18], activateOut_17r, activateOut_17a);
  selem I20 (sreq_0n[16], sreq_0n[17], activateOut_16r, activateOut_16a);
  selem I21 (sreq_0n[15], sreq_0n[16], activateOut_15r, activateOut_15a);
  selem I22 (sreq_0n[14], sreq_0n[15], activateOut_14r, activateOut_14a);
  selem I23 (sreq_0n[13], sreq_0n[14], activateOut_13r, activateOut_13a);
  selem I24 (sreq_0n[12], sreq_0n[13], activateOut_12r, activateOut_12a);
  selem I25 (sreq_0n[11], sreq_0n[12], activateOut_11r, activateOut_11a);
  selem I26 (sreq_0n[10], sreq_0n[11], activateOut_10r, activateOut_10a);
  selem I27 (sreq_0n[9], sreq_0n[10], activateOut_9r, activateOut_9a);
  selem I28 (sreq_0n[8], sreq_0n[9], activateOut_8r, activateOut_8a);
  selem I29 (sreq_0n[7], sreq_0n[8], activateOut_7r, activateOut_7a);
  selem I30 (sreq_0n[6], sreq_0n[7], activateOut_6r, activateOut_6a);
  selem I31 (sreq_0n[5], sreq_0n[6], activateOut_5r, activateOut_5a);
  selem I32 (sreq_0n[4], sreq_0n[5], activateOut_4r, activateOut_4a);
  selem I33 (sreq_0n[3], sreq_0n[4], activateOut_3r, activateOut_3a);
  selem I34 (sreq_0n[2], sreq_0n[3], activateOut_2r, activateOut_2a);
  selem I35 (sreq_0n[1], sreq_0n[2], activateOut_1r, activateOut_1a);
  selem I36 (sreq_0n[0], sreq_0n[1], activateOut_0r, activateOut_0a);
endmodule

module BrzSlice_1_34_32 (
  out_0r, out_0a, out_0d,
  inp_0r, inp_0a, inp_0d
);
  input out_0r;
  output out_0a;
  output out_0d;
  output inp_0r;
  input inp_0a;
  input [33:0] inp_0d;
  assign inp_0r = out_0r;
  assign out_0a = inp_0a;
  assign out_0d = inp_0d[32];
endmodule

module BrzSlice_32_34_1 (
  out_0r, out_0a, out_0d,
  inp_0r, inp_0a, inp_0d
);
  input out_0r;
  output out_0a;
  output [31:0] out_0d;
  output inp_0r;
  input inp_0a;
  input [33:0] inp_0d;
  assign inp_0r = out_0r;
  assign out_0a = inp_0a;
  assign out_0d[0] = inp_0d[1];
  assign out_0d[1] = inp_0d[2];
  assign out_0d[2] = inp_0d[3];
  assign out_0d[3] = inp_0d[4];
  assign out_0d[4] = inp_0d[5];
  assign out_0d[5] = inp_0d[6];
  assign out_0d[6] = inp_0d[7];
  assign out_0d[7] = inp_0d[8];
  assign out_0d[8] = inp_0d[9];
  assign out_0d[9] = inp_0d[10];
  assign out_0d[10] = inp_0d[11];
  assign out_0d[11] = inp_0d[12];
  assign out_0d[12] = inp_0d[13];
  assign out_0d[13] = inp_0d[14];
  assign out_0d[14] = inp_0d[15];
  assign out_0d[15] = inp_0d[16];
  assign out_0d[16] = inp_0d[17];
  assign out_0d[17] = inp_0d[18];
  assign out_0d[18] = inp_0d[19];
  assign out_0d[19] = inp_0d[20];
  assign out_0d[20] = inp_0d[21];
  assign out_0d[21] = inp_0d[22];
  assign out_0d[22] = inp_0d[23];
  assign out_0d[23] = inp_0d[24];
  assign out_0d[24] = inp_0d[25];
  assign out_0d[25] = inp_0d[26];
  assign out_0d[26] = inp_0d[27];
  assign out_0d[27] = inp_0d[28];
  assign out_0d[28] = inp_0d[29];
  assign out_0d[29] = inp_0d[30];
  assign out_0d[30] = inp_0d[31];
  assign out_0d[31] = inp_0d[32];
endmodule

module BrzUnaryFunc_1_1_s6_Invert_s5_false (
  out_0r, out_0a, out_0d,
  inp_0r, inp_0a, inp_0d
);
  input out_0r;
  output out_0a;
  output out_0d;
  output inp_0r;
  input inp_0a;
  input inp_0d;
  wire nStart_0n;
  wire [1:0] nCv_0n;
  wire [1:0] c_0n;
  wire i_0n;
  wire j_0n;
  wire start_0n;
  wire done_0n;
  IV I0 (out_0d, inp_0d);
  assign done_0n = start_0n;
  assign out_0a = done_0n;
  assign start_0n = inp_0a;
  assign inp_0r = out_0r;
endmodule

module BrzUnaryFunc_16_16_s6_Negate_s4_true (
  out_0r, out_0a, out_0d,
  inp_0r, inp_0a, inp_0d
);
  input out_0r;
  output out_0a;
  output [15:0] out_0d;
  output inp_0r;
  input inp_0a;
  input [15:0] inp_0d;
  wire [3:0] internal_0n;
  wire nStart_0n;
  wire [16:0] nCv_0n;
  wire [16:0] c_0n;
  wire [15:0] i_0n;
  wire [15:0] j_0n;
  wire start_0n;
  wire done_0n;
  wire gnd;
  wire vcc;
  GND gnd_cell_instance (gnd);
  VCC vcc_cell_instance (vcc);
  NR4 I0 (internal_0n[0], nCv_0n[1], nCv_0n[2], nCv_0n[3], nCv_0n[4]);
  NR4 I1 (internal_0n[1], nCv_0n[5], nCv_0n[6], nCv_0n[7], nCv_0n[8]);
  NR4 I2 (internal_0n[2], nCv_0n[9], nCv_0n[10], nCv_0n[11], nCv_0n[12]);
  NR4 I3 (internal_0n[3], nCv_0n[13], nCv_0n[14], nCv_0n[15], nCv_0n[16]);
  AN4 I4 (done_0n, internal_0n[0], internal_0n[1], internal_0n[2], internal_0n[3]);
  balsa_fa I5 (nStart_0n, i_0n[0], j_0n[0], nCv_0n[0], c_0n[0], nCv_0n[1], c_0n[1], out_0d[0]);
  balsa_fa I6 (nStart_0n, i_0n[1], j_0n[1], nCv_0n[1], c_0n[1], nCv_0n[2], c_0n[2], out_0d[1]);
  balsa_fa I7 (nStart_0n, i_0n[2], j_0n[2], nCv_0n[2], c_0n[2], nCv_0n[3], c_0n[3], out_0d[2]);
  balsa_fa I8 (nStart_0n, i_0n[3], j_0n[3], nCv_0n[3], c_0n[3], nCv_0n[4], c_0n[4], out_0d[3]);
  balsa_fa I9 (nStart_0n, i_0n[4], j_0n[4], nCv_0n[4], c_0n[4], nCv_0n[5], c_0n[5], out_0d[4]);
  balsa_fa I10 (nStart_0n, i_0n[5], j_0n[5], nCv_0n[5], c_0n[5], nCv_0n[6], c_0n[6], out_0d[5]);
  balsa_fa I11 (nStart_0n, i_0n[6], j_0n[6], nCv_0n[6], c_0n[6], nCv_0n[7], c_0n[7], out_0d[6]);
  balsa_fa I12 (nStart_0n, i_0n[7], j_0n[7], nCv_0n[7], c_0n[7], nCv_0n[8], c_0n[8], out_0d[7]);
  balsa_fa I13 (nStart_0n, i_0n[8], j_0n[8], nCv_0n[8], c_0n[8], nCv_0n[9], c_0n[9], out_0d[8]);
  balsa_fa I14 (nStart_0n, i_0n[9], j_0n[9], nCv_0n[9], c_0n[9], nCv_0n[10], c_0n[10], out_0d[9]);
  balsa_fa I15 (nStart_0n, i_0n[10], j_0n[10], nCv_0n[10], c_0n[10], nCv_0n[11], c_0n[11], out_0d[10]);
  balsa_fa I16 (nStart_0n, i_0n[11], j_0n[11], nCv_0n[11], c_0n[11], nCv_0n[12], c_0n[12], out_0d[11]);
  balsa_fa I17 (nStart_0n, i_0n[12], j_0n[12], nCv_0n[12], c_0n[12], nCv_0n[13], c_0n[13], out_0d[12]);
  balsa_fa I18 (nStart_0n, i_0n[13], j_0n[13], nCv_0n[13], c_0n[13], nCv_0n[14], c_0n[14], out_0d[13]);
  balsa_fa I19 (nStart_0n, i_0n[14], j_0n[14], nCv_0n[14], c_0n[14], nCv_0n[15], c_0n[15], out_0d[14]);
  balsa_fa I20 (nStart_0n, i_0n[15], j_0n[15], nCv_0n[15], c_0n[15], nCv_0n[16], c_0n[16], out_0d[15]);
  assign c_0n[0] = vcc;
  assign j_0n[0] = gnd;
  assign j_0n[1] = gnd;
  assign j_0n[2] = gnd;
  assign j_0n[3] = gnd;
  assign j_0n[4] = gnd;
  assign j_0n[5] = gnd;
  assign j_0n[6] = gnd;
  assign j_0n[7] = gnd;
  assign j_0n[8] = gnd;
  assign j_0n[9] = gnd;
  assign j_0n[10] = gnd;
  assign j_0n[11] = gnd;
  assign j_0n[12] = gnd;
  assign j_0n[13] = gnd;
  assign j_0n[14] = gnd;
  assign j_0n[15] = gnd;
  assign nCv_0n[0] = nStart_0n;
  IV I39 (i_0n[0], inp_0d[0]);
  IV I40 (i_0n[1], inp_0d[1]);
  IV I41 (i_0n[2], inp_0d[2]);
  IV I42 (i_0n[3], inp_0d[3]);
  IV I43 (i_0n[4], inp_0d[4]);
  IV I44 (i_0n[5], inp_0d[5]);
  IV I45 (i_0n[6], inp_0d[6]);
  IV I46 (i_0n[7], inp_0d[7]);
  IV I47 (i_0n[8], inp_0d[8]);
  IV I48 (i_0n[9], inp_0d[9]);
  IV I49 (i_0n[10], inp_0d[10]);
  IV I50 (i_0n[11], inp_0d[11]);
  IV I51 (i_0n[12], inp_0d[12]);
  IV I52 (i_0n[13], inp_0d[13]);
  IV I53 (i_0n[14], inp_0d[14]);
  IV I54 (i_0n[15], inp_0d[15]);
  IV I55 (nStart_0n, start_0n);
  assign out_0a = done_0n;
  assign start_0n = inp_0a;
  assign inp_0r = out_0r;
endmodule

module BrzVariable_1_1_s0_ (
  write_0r, write_0a, write_0d,
  read_0r, read_0a, read_0d
);
  input write_0r;
  output write_0a;
  input write_0d;
  input read_0r;
  output read_0a;
  output read_0d;
  wire data_0n;
  wire nWriteReq_0n;
  wire bWriteReq_0n;
  wire nbWriteReq_0n;
  assign read_0a = read_0r;
  assign read_0d = data_0n;
  LD1 I2 (write_0d, bWriteReq_0n, data_0n);
  IV I3 (write_0a, nbWriteReq_0n);
  IV I4 (nbWriteReq_0n, bWriteReq_0n);
  IV I5 (bWriteReq_0n, nWriteReq_0n);
  IV I6 (nWriteReq_0n, write_0r);
endmodule

module BrzVariable_16_1_s0_ (
  write_0r, write_0a, write_0d,
  read_0r, read_0a, read_0d
);
  input write_0r;
  output write_0a;
  input [15:0] write_0d;
  input read_0r;
  output read_0a;
  output [15:0] read_0d;
  wire [15:0] data_0n;
  wire nWriteReq_0n;
  wire bWriteReq_0n;
  wire nbWriteReq_0n;
  assign read_0a = read_0r;
  assign read_0d[0] = data_0n[0];
  assign read_0d[1] = data_0n[1];
  assign read_0d[2] = data_0n[2];
  assign read_0d[3] = data_0n[3];
  assign read_0d[4] = data_0n[4];
  assign read_0d[5] = data_0n[5];
  assign read_0d[6] = data_0n[6];
  assign read_0d[7] = data_0n[7];
  assign read_0d[8] = data_0n[8];
  assign read_0d[9] = data_0n[9];
  assign read_0d[10] = data_0n[10];
  assign read_0d[11] = data_0n[11];
  assign read_0d[12] = data_0n[12];
  assign read_0d[13] = data_0n[13];
  assign read_0d[14] = data_0n[14];
  assign read_0d[15] = data_0n[15];
  LD1 I17 (write_0d[0], bWriteReq_0n, data_0n[0]);
  LD1 I18 (write_0d[1], bWriteReq_0n, data_0n[1]);
  LD1 I19 (write_0d[2], bWriteReq_0n, data_0n[2]);
  LD1 I20 (write_0d[3], bWriteReq_0n, data_0n[3]);
  LD1 I21 (write_0d[4], bWriteReq_0n, data_0n[4]);
  LD1 I22 (write_0d[5], bWriteReq_0n, data_0n[5]);
  LD1 I23 (write_0d[6], bWriteReq_0n, data_0n[6]);
  LD1 I24 (write_0d[7], bWriteReq_0n, data_0n[7]);
  LD1 I25 (write_0d[8], bWriteReq_0n, data_0n[8]);
  LD1 I26 (write_0d[9], bWriteReq_0n, data_0n[9]);
  LD1 I27 (write_0d[10], bWriteReq_0n, data_0n[10]);
  LD1 I28 (write_0d[11], bWriteReq_0n, data_0n[11]);
  LD1 I29 (write_0d[12], bWriteReq_0n, data_0n[12]);
  LD1 I30 (write_0d[13], bWriteReq_0n, data_0n[13]);
  LD1 I31 (write_0d[14], bWriteReq_0n, data_0n[14]);
  LD1 I32 (write_0d[15], bWriteReq_0n, data_0n[15]);
  IV I33 (write_0a, nbWriteReq_0n);
  IV I34 (nbWriteReq_0n, bWriteReq_0n);
  IV I35 (bWriteReq_0n, nWriteReq_0n);
  IV I36 (nWriteReq_0n, write_0r);
endmodule

module BrzVariable_16_2_s0_ (
  write_0r, write_0a, write_0d,
  read_0r, read_0a, read_0d,
  read_1r, read_1a, read_1d
);
  input write_0r;
  output write_0a;
  input [15:0] write_0d;
  input read_0r;
  output read_0a;
  output [15:0] read_0d;
  input read_1r;
  output read_1a;
  output [15:0] read_1d;
  wire [15:0] data_0n;
  wire nWriteReq_0n;
  wire bWriteReq_0n;
  wire nbWriteReq_0n;
  assign read_0a = read_0r;
  assign read_1a = read_1r;
  assign read_1d[0] = data_0n[0];
  assign read_1d[1] = data_0n[1];
  assign read_1d[2] = data_0n[2];
  assign read_1d[3] = data_0n[3];
  assign read_1d[4] = data_0n[4];
  assign read_1d[5] = data_0n[5];
  assign read_1d[6] = data_0n[6];
  assign read_1d[7] = data_0n[7];
  assign read_1d[8] = data_0n[8];
  assign read_1d[9] = data_0n[9];
  assign read_1d[10] = data_0n[10];
  assign read_1d[11] = data_0n[11];
  assign read_1d[12] = data_0n[12];
  assign read_1d[13] = data_0n[13];
  assign read_1d[14] = data_0n[14];
  assign read_1d[15] = data_0n[15];
  assign read_0d[0] = data_0n[0];
  assign read_0d[1] = data_0n[1];
  assign read_0d[2] = data_0n[2];
  assign read_0d[3] = data_0n[3];
  assign read_0d[4] = data_0n[4];
  assign read_0d[5] = data_0n[5];
  assign read_0d[6] = data_0n[6];
  assign read_0d[7] = data_0n[7];
  assign read_0d[8] = data_0n[8];
  assign read_0d[9] = data_0n[9];
  assign read_0d[10] = data_0n[10];
  assign read_0d[11] = data_0n[11];
  assign read_0d[12] = data_0n[12];
  assign read_0d[13] = data_0n[13];
  assign read_0d[14] = data_0n[14];
  assign read_0d[15] = data_0n[15];
  LD1 I34 (write_0d[0], bWriteReq_0n, data_0n[0]);
  LD1 I35 (write_0d[1], bWriteReq_0n, data_0n[1]);
  LD1 I36 (write_0d[2], bWriteReq_0n, data_0n[2]);
  LD1 I37 (write_0d[3], bWriteReq_0n, data_0n[3]);
  LD1 I38 (write_0d[4], bWriteReq_0n, data_0n[4]);
  LD1 I39 (write_0d[5], bWriteReq_0n, data_0n[5]);
  LD1 I40 (write_0d[6], bWriteReq_0n, data_0n[6]);
  LD1 I41 (write_0d[7], bWriteReq_0n, data_0n[7]);
  LD1 I42 (write_0d[8], bWriteReq_0n, data_0n[8]);
  LD1 I43 (write_0d[9], bWriteReq_0n, data_0n[9]);
  LD1 I44 (write_0d[10], bWriteReq_0n, data_0n[10]);
  LD1 I45 (write_0d[11], bWriteReq_0n, data_0n[11]);
  LD1 I46 (write_0d[12], bWriteReq_0n, data_0n[12]);
  LD1 I47 (write_0d[13], bWriteReq_0n, data_0n[13]);
  LD1 I48 (write_0d[14], bWriteReq_0n, data_0n[14]);
  LD1 I49 (write_0d[15], bWriteReq_0n, data_0n[15]);
  IV I50 (write_0a, nbWriteReq_0n);
  IV I51 (nbWriteReq_0n, bWriteReq_0n);
  IV I52 (bWriteReq_0n, nWriteReq_0n);
  IV I53 (nWriteReq_0n, write_0r);
endmodule

module BrzVariable_33_1_s0_ (
  write_0r, write_0a, write_0d,
  read_0r, read_0a, read_0d
);
  input write_0r;
  output write_0a;
  input [32:0] write_0d;
  input read_0r;
  output read_0a;
  output [32:0] read_0d;
  wire [32:0] data_0n;
  wire nWriteReq_0n;
  wire bWriteReq_0n;
  wire nbWriteReq_0n;
  assign read_0a = read_0r;
  assign read_0d[0] = data_0n[0];
  assign read_0d[1] = data_0n[1];
  assign read_0d[2] = data_0n[2];
  assign read_0d[3] = data_0n[3];
  assign read_0d[4] = data_0n[4];
  assign read_0d[5] = data_0n[5];
  assign read_0d[6] = data_0n[6];
  assign read_0d[7] = data_0n[7];
  assign read_0d[8] = data_0n[8];
  assign read_0d[9] = data_0n[9];
  assign read_0d[10] = data_0n[10];
  assign read_0d[11] = data_0n[11];
  assign read_0d[12] = data_0n[12];
  assign read_0d[13] = data_0n[13];
  assign read_0d[14] = data_0n[14];
  assign read_0d[15] = data_0n[15];
  assign read_0d[16] = data_0n[16];
  assign read_0d[17] = data_0n[17];
  assign read_0d[18] = data_0n[18];
  assign read_0d[19] = data_0n[19];
  assign read_0d[20] = data_0n[20];
  assign read_0d[21] = data_0n[21];
  assign read_0d[22] = data_0n[22];
  assign read_0d[23] = data_0n[23];
  assign read_0d[24] = data_0n[24];
  assign read_0d[25] = data_0n[25];
  assign read_0d[26] = data_0n[26];
  assign read_0d[27] = data_0n[27];
  assign read_0d[28] = data_0n[28];
  assign read_0d[29] = data_0n[29];
  assign read_0d[30] = data_0n[30];
  assign read_0d[31] = data_0n[31];
  assign read_0d[32] = data_0n[32];
  LD1 I34 (write_0d[0], bWriteReq_0n, data_0n[0]);
  LD1 I35 (write_0d[1], bWriteReq_0n, data_0n[1]);
  LD1 I36 (write_0d[2], bWriteReq_0n, data_0n[2]);
  LD1 I37 (write_0d[3], bWriteReq_0n, data_0n[3]);
  LD1 I38 (write_0d[4], bWriteReq_0n, data_0n[4]);
  LD1 I39 (write_0d[5], bWriteReq_0n, data_0n[5]);
  LD1 I40 (write_0d[6], bWriteReq_0n, data_0n[6]);
  LD1 I41 (write_0d[7], bWriteReq_0n, data_0n[7]);
  LD1 I42 (write_0d[8], bWriteReq_0n, data_0n[8]);
  LD1 I43 (write_0d[9], bWriteReq_0n, data_0n[9]);
  LD1 I44 (write_0d[10], bWriteReq_0n, data_0n[10]);
  LD1 I45 (write_0d[11], bWriteReq_0n, data_0n[11]);
  LD1 I46 (write_0d[12], bWriteReq_0n, data_0n[12]);
  LD1 I47 (write_0d[13], bWriteReq_0n, data_0n[13]);
  LD1 I48 (write_0d[14], bWriteReq_0n, data_0n[14]);
  LD1 I49 (write_0d[15], bWriteReq_0n, data_0n[15]);
  LD1 I50 (write_0d[16], bWriteReq_0n, data_0n[16]);
  LD1 I51 (write_0d[17], bWriteReq_0n, data_0n[17]);
  LD1 I52 (write_0d[18], bWriteReq_0n, data_0n[18]);
  LD1 I53 (write_0d[19], bWriteReq_0n, data_0n[19]);
  LD1 I54 (write_0d[20], bWriteReq_0n, data_0n[20]);
  LD1 I55 (write_0d[21], bWriteReq_0n, data_0n[21]);
  LD1 I56 (write_0d[22], bWriteReq_0n, data_0n[22]);
  LD1 I57 (write_0d[23], bWriteReq_0n, data_0n[23]);
  LD1 I58 (write_0d[24], bWriteReq_0n, data_0n[24]);
  LD1 I59 (write_0d[25], bWriteReq_0n, data_0n[25]);
  LD1 I60 (write_0d[26], bWriteReq_0n, data_0n[26]);
  LD1 I61 (write_0d[27], bWriteReq_0n, data_0n[27]);
  LD1 I62 (write_0d[28], bWriteReq_0n, data_0n[28]);
  LD1 I63 (write_0d[29], bWriteReq_0n, data_0n[29]);
  LD1 I64 (write_0d[30], bWriteReq_0n, data_0n[30]);
  LD1 I65 (write_0d[31], bWriteReq_0n, data_0n[31]);
  LD1 I66 (write_0d[32], bWriteReq_0n, data_0n[32]);
  IV I67 (write_0a, nbWriteReq_0n);
  IV I68 (nbWriteReq_0n, bWriteReq_0n);
  IV I69 (bWriteReq_0n, nWriteReq_0n);
  IV I70 (nWriteReq_0n, write_0r);
endmodule

module BrzVariable_33_32_s0_ (
  write_0r, write_0a, write_0d,
  read_0r, read_0a, read_0d,
  read_1r, read_1a, read_1d,
  read_2r, read_2a, read_2d,
  read_3r, read_3a, read_3d,
  read_4r, read_4a, read_4d,
  read_5r, read_5a, read_5d,
  read_6r, read_6a, read_6d,
  read_7r, read_7a, read_7d,
  read_8r, read_8a, read_8d,
  read_9r, read_9a, read_9d,
  read_10r, read_10a, read_10d,
  read_11r, read_11a, read_11d,
  read_12r, read_12a, read_12d,
  read_13r, read_13a, read_13d,
  read_14r, read_14a, read_14d,
  read_15r, read_15a, read_15d,
  read_16r, read_16a, read_16d,
  read_17r, read_17a, read_17d,
  read_18r, read_18a, read_18d,
  read_19r, read_19a, read_19d,
  read_20r, read_20a, read_20d,
  read_21r, read_21a, read_21d,
  read_22r, read_22a, read_22d,
  read_23r, read_23a, read_23d,
  read_24r, read_24a, read_24d,
  read_25r, read_25a, read_25d,
  read_26r, read_26a, read_26d,
  read_27r, read_27a, read_27d,
  read_28r, read_28a, read_28d,
  read_29r, read_29a, read_29d,
  read_30r, read_30a, read_30d,
  read_31r, read_31a, read_31d
);
  input write_0r;
  output write_0a;
  input [32:0] write_0d;
  input read_0r;
  output read_0a;
  output [32:0] read_0d;
  input read_1r;
  output read_1a;
  output [32:0] read_1d;
  input read_2r;
  output read_2a;
  output [32:0] read_2d;
  input read_3r;
  output read_3a;
  output [32:0] read_3d;
  input read_4r;
  output read_4a;
  output [32:0] read_4d;
  input read_5r;
  output read_5a;
  output [32:0] read_5d;
  input read_6r;
  output read_6a;
  output [32:0] read_6d;
  input read_7r;
  output read_7a;
  output [32:0] read_7d;
  input read_8r;
  output read_8a;
  output [32:0] read_8d;
  input read_9r;
  output read_9a;
  output [32:0] read_9d;
  input read_10r;
  output read_10a;
  output [32:0] read_10d;
  input read_11r;
  output read_11a;
  output [32:0] read_11d;
  input read_12r;
  output read_12a;
  output [32:0] read_12d;
  input read_13r;
  output read_13a;
  output [32:0] read_13d;
  input read_14r;
  output read_14a;
  output [32:0] read_14d;
  input read_15r;
  output read_15a;
  output [32:0] read_15d;
  input read_16r;
  output read_16a;
  output [32:0] read_16d;
  input read_17r;
  output read_17a;
  output [32:0] read_17d;
  input read_18r;
  output read_18a;
  output [32:0] read_18d;
  input read_19r;
  output read_19a;
  output [32:0] read_19d;
  input read_20r;
  output read_20a;
  output [32:0] read_20d;
  input read_21r;
  output read_21a;
  output [32:0] read_21d;
  input read_22r;
  output read_22a;
  output [32:0] read_22d;
  input read_23r;
  output read_23a;
  output [32:0] read_23d;
  input read_24r;
  output read_24a;
  output [32:0] read_24d;
  input read_25r;
  output read_25a;
  output [32:0] read_25d;
  input read_26r;
  output read_26a;
  output [32:0] read_26d;
  input read_27r;
  output read_27a;
  output [32:0] read_27d;
  input read_28r;
  output read_28a;
  output [32:0] read_28d;
  input read_29r;
  output read_29a;
  output [32:0] read_29d;
  input read_30r;
  output read_30a;
  output [32:0] read_30d;
  input read_31r;
  output read_31a;
  output [32:0] read_31d;
  wire [32:0] data_0n;
  wire nWriteReq_0n;
  wire bWriteReq_0n;
  wire nbWriteReq_0n;
  assign read_0a = read_0r;
  assign read_1a = read_1r;
  assign read_2a = read_2r;
  assign read_3a = read_3r;
  assign read_4a = read_4r;
  assign read_5a = read_5r;
  assign read_6a = read_6r;
  assign read_7a = read_7r;
  assign read_8a = read_8r;
  assign read_9a = read_9r;
  assign read_10a = read_10r;
  assign read_11a = read_11r;
  assign read_12a = read_12r;
  assign read_13a = read_13r;
  assign read_14a = read_14r;
  assign read_15a = read_15r;
  assign read_16a = read_16r;
  assign read_17a = read_17r;
  assign read_18a = read_18r;
  assign read_19a = read_19r;
  assign read_20a = read_20r;
  assign read_21a = read_21r;
  assign read_22a = read_22r;
  assign read_23a = read_23r;
  assign read_24a = read_24r;
  assign read_25a = read_25r;
  assign read_26a = read_26r;
  assign read_27a = read_27r;
  assign read_28a = read_28r;
  assign read_29a = read_29r;
  assign read_30a = read_30r;
  assign read_31a = read_31r;
  assign read_31d[0] = data_0n[0];
  assign read_31d[1] = data_0n[1];
  assign read_31d[2] = data_0n[2];
  assign read_31d[3] = data_0n[3];
  assign read_31d[4] = data_0n[4];
  assign read_31d[5] = data_0n[5];
  assign read_31d[6] = data_0n[6];
  assign read_31d[7] = data_0n[7];
  assign read_31d[8] = data_0n[8];
  assign read_31d[9] = data_0n[9];
  assign read_31d[10] = data_0n[10];
  assign read_31d[11] = data_0n[11];
  assign read_31d[12] = data_0n[12];
  assign read_31d[13] = data_0n[13];
  assign read_31d[14] = data_0n[14];
  assign read_31d[15] = data_0n[15];
  assign read_31d[16] = data_0n[16];
  assign read_31d[17] = data_0n[17];
  assign read_31d[18] = data_0n[18];
  assign read_31d[19] = data_0n[19];
  assign read_31d[20] = data_0n[20];
  assign read_31d[21] = data_0n[21];
  assign read_31d[22] = data_0n[22];
  assign read_31d[23] = data_0n[23];
  assign read_31d[24] = data_0n[24];
  assign read_31d[25] = data_0n[25];
  assign read_31d[26] = data_0n[26];
  assign read_31d[27] = data_0n[27];
  assign read_31d[28] = data_0n[28];
  assign read_31d[29] = data_0n[29];
  assign read_31d[30] = data_0n[30];
  assign read_31d[31] = data_0n[31];
  assign read_31d[32] = data_0n[32];
  assign read_30d[0] = data_0n[0];
  assign read_30d[1] = data_0n[1];
  assign read_30d[2] = data_0n[2];
  assign read_30d[3] = data_0n[3];
  assign read_30d[4] = data_0n[4];
  assign read_30d[5] = data_0n[5];
  assign read_30d[6] = data_0n[6];
  assign read_30d[7] = data_0n[7];
  assign read_30d[8] = data_0n[8];
  assign read_30d[9] = data_0n[9];
  assign read_30d[10] = data_0n[10];
  assign read_30d[11] = data_0n[11];
  assign read_30d[12] = data_0n[12];
  assign read_30d[13] = data_0n[13];
  assign read_30d[14] = data_0n[14];
  assign read_30d[15] = data_0n[15];
  assign read_30d[16] = data_0n[16];
  assign read_30d[17] = data_0n[17];
  assign read_30d[18] = data_0n[18];
  assign read_30d[19] = data_0n[19];
  assign read_30d[20] = data_0n[20];
  assign read_30d[21] = data_0n[21];
  assign read_30d[22] = data_0n[22];
  assign read_30d[23] = data_0n[23];
  assign read_30d[24] = data_0n[24];
  assign read_30d[25] = data_0n[25];
  assign read_30d[26] = data_0n[26];
  assign read_30d[27] = data_0n[27];
  assign read_30d[28] = data_0n[28];
  assign read_30d[29] = data_0n[29];
  assign read_30d[30] = data_0n[30];
  assign read_30d[31] = data_0n[31];
  assign read_30d[32] = data_0n[32];
  assign read_29d[0] = data_0n[0];
  assign read_29d[1] = data_0n[1];
  assign read_29d[2] = data_0n[2];
  assign read_29d[3] = data_0n[3];
  assign read_29d[4] = data_0n[4];
  assign read_29d[5] = data_0n[5];
  assign read_29d[6] = data_0n[6];
  assign read_29d[7] = data_0n[7];
  assign read_29d[8] = data_0n[8];
  assign read_29d[9] = data_0n[9];
  assign read_29d[10] = data_0n[10];
  assign read_29d[11] = data_0n[11];
  assign read_29d[12] = data_0n[12];
  assign read_29d[13] = data_0n[13];
  assign read_29d[14] = data_0n[14];
  assign read_29d[15] = data_0n[15];
  assign read_29d[16] = data_0n[16];
  assign read_29d[17] = data_0n[17];
  assign read_29d[18] = data_0n[18];
  assign read_29d[19] = data_0n[19];
  assign read_29d[20] = data_0n[20];
  assign read_29d[21] = data_0n[21];
  assign read_29d[22] = data_0n[22];
  assign read_29d[23] = data_0n[23];
  assign read_29d[24] = data_0n[24];
  assign read_29d[25] = data_0n[25];
  assign read_29d[26] = data_0n[26];
  assign read_29d[27] = data_0n[27];
  assign read_29d[28] = data_0n[28];
  assign read_29d[29] = data_0n[29];
  assign read_29d[30] = data_0n[30];
  assign read_29d[31] = data_0n[31];
  assign read_29d[32] = data_0n[32];
  assign read_28d[0] = data_0n[0];
  assign read_28d[1] = data_0n[1];
  assign read_28d[2] = data_0n[2];
  assign read_28d[3] = data_0n[3];
  assign read_28d[4] = data_0n[4];
  assign read_28d[5] = data_0n[5];
  assign read_28d[6] = data_0n[6];
  assign read_28d[7] = data_0n[7];
  assign read_28d[8] = data_0n[8];
  assign read_28d[9] = data_0n[9];
  assign read_28d[10] = data_0n[10];
  assign read_28d[11] = data_0n[11];
  assign read_28d[12] = data_0n[12];
  assign read_28d[13] = data_0n[13];
  assign read_28d[14] = data_0n[14];
  assign read_28d[15] = data_0n[15];
  assign read_28d[16] = data_0n[16];
  assign read_28d[17] = data_0n[17];
  assign read_28d[18] = data_0n[18];
  assign read_28d[19] = data_0n[19];
  assign read_28d[20] = data_0n[20];
  assign read_28d[21] = data_0n[21];
  assign read_28d[22] = data_0n[22];
  assign read_28d[23] = data_0n[23];
  assign read_28d[24] = data_0n[24];
  assign read_28d[25] = data_0n[25];
  assign read_28d[26] = data_0n[26];
  assign read_28d[27] = data_0n[27];
  assign read_28d[28] = data_0n[28];
  assign read_28d[29] = data_0n[29];
  assign read_28d[30] = data_0n[30];
  assign read_28d[31] = data_0n[31];
  assign read_28d[32] = data_0n[32];
  assign read_27d[0] = data_0n[0];
  assign read_27d[1] = data_0n[1];
  assign read_27d[2] = data_0n[2];
  assign read_27d[3] = data_0n[3];
  assign read_27d[4] = data_0n[4];
  assign read_27d[5] = data_0n[5];
  assign read_27d[6] = data_0n[6];
  assign read_27d[7] = data_0n[7];
  assign read_27d[8] = data_0n[8];
  assign read_27d[9] = data_0n[9];
  assign read_27d[10] = data_0n[10];
  assign read_27d[11] = data_0n[11];
  assign read_27d[12] = data_0n[12];
  assign read_27d[13] = data_0n[13];
  assign read_27d[14] = data_0n[14];
  assign read_27d[15] = data_0n[15];
  assign read_27d[16] = data_0n[16];
  assign read_27d[17] = data_0n[17];
  assign read_27d[18] = data_0n[18];
  assign read_27d[19] = data_0n[19];
  assign read_27d[20] = data_0n[20];
  assign read_27d[21] = data_0n[21];
  assign read_27d[22] = data_0n[22];
  assign read_27d[23] = data_0n[23];
  assign read_27d[24] = data_0n[24];
  assign read_27d[25] = data_0n[25];
  assign read_27d[26] = data_0n[26];
  assign read_27d[27] = data_0n[27];
  assign read_27d[28] = data_0n[28];
  assign read_27d[29] = data_0n[29];
  assign read_27d[30] = data_0n[30];
  assign read_27d[31] = data_0n[31];
  assign read_27d[32] = data_0n[32];
  assign read_26d[0] = data_0n[0];
  assign read_26d[1] = data_0n[1];
  assign read_26d[2] = data_0n[2];
  assign read_26d[3] = data_0n[3];
  assign read_26d[4] = data_0n[4];
  assign read_26d[5] = data_0n[5];
  assign read_26d[6] = data_0n[6];
  assign read_26d[7] = data_0n[7];
  assign read_26d[8] = data_0n[8];
  assign read_26d[9] = data_0n[9];
  assign read_26d[10] = data_0n[10];
  assign read_26d[11] = data_0n[11];
  assign read_26d[12] = data_0n[12];
  assign read_26d[13] = data_0n[13];
  assign read_26d[14] = data_0n[14];
  assign read_26d[15] = data_0n[15];
  assign read_26d[16] = data_0n[16];
  assign read_26d[17] = data_0n[17];
  assign read_26d[18] = data_0n[18];
  assign read_26d[19] = data_0n[19];
  assign read_26d[20] = data_0n[20];
  assign read_26d[21] = data_0n[21];
  assign read_26d[22] = data_0n[22];
  assign read_26d[23] = data_0n[23];
  assign read_26d[24] = data_0n[24];
  assign read_26d[25] = data_0n[25];
  assign read_26d[26] = data_0n[26];
  assign read_26d[27] = data_0n[27];
  assign read_26d[28] = data_0n[28];
  assign read_26d[29] = data_0n[29];
  assign read_26d[30] = data_0n[30];
  assign read_26d[31] = data_0n[31];
  assign read_26d[32] = data_0n[32];
  assign read_25d[0] = data_0n[0];
  assign read_25d[1] = data_0n[1];
  assign read_25d[2] = data_0n[2];
  assign read_25d[3] = data_0n[3];
  assign read_25d[4] = data_0n[4];
  assign read_25d[5] = data_0n[5];
  assign read_25d[6] = data_0n[6];
  assign read_25d[7] = data_0n[7];
  assign read_25d[8] = data_0n[8];
  assign read_25d[9] = data_0n[9];
  assign read_25d[10] = data_0n[10];
  assign read_25d[11] = data_0n[11];
  assign read_25d[12] = data_0n[12];
  assign read_25d[13] = data_0n[13];
  assign read_25d[14] = data_0n[14];
  assign read_25d[15] = data_0n[15];
  assign read_25d[16] = data_0n[16];
  assign read_25d[17] = data_0n[17];
  assign read_25d[18] = data_0n[18];
  assign read_25d[19] = data_0n[19];
  assign read_25d[20] = data_0n[20];
  assign read_25d[21] = data_0n[21];
  assign read_25d[22] = data_0n[22];
  assign read_25d[23] = data_0n[23];
  assign read_25d[24] = data_0n[24];
  assign read_25d[25] = data_0n[25];
  assign read_25d[26] = data_0n[26];
  assign read_25d[27] = data_0n[27];
  assign read_25d[28] = data_0n[28];
  assign read_25d[29] = data_0n[29];
  assign read_25d[30] = data_0n[30];
  assign read_25d[31] = data_0n[31];
  assign read_25d[32] = data_0n[32];
  assign read_24d[0] = data_0n[0];
  assign read_24d[1] = data_0n[1];
  assign read_24d[2] = data_0n[2];
  assign read_24d[3] = data_0n[3];
  assign read_24d[4] = data_0n[4];
  assign read_24d[5] = data_0n[5];
  assign read_24d[6] = data_0n[6];
  assign read_24d[7] = data_0n[7];
  assign read_24d[8] = data_0n[8];
  assign read_24d[9] = data_0n[9];
  assign read_24d[10] = data_0n[10];
  assign read_24d[11] = data_0n[11];
  assign read_24d[12] = data_0n[12];
  assign read_24d[13] = data_0n[13];
  assign read_24d[14] = data_0n[14];
  assign read_24d[15] = data_0n[15];
  assign read_24d[16] = data_0n[16];
  assign read_24d[17] = data_0n[17];
  assign read_24d[18] = data_0n[18];
  assign read_24d[19] = data_0n[19];
  assign read_24d[20] = data_0n[20];
  assign read_24d[21] = data_0n[21];
  assign read_24d[22] = data_0n[22];
  assign read_24d[23] = data_0n[23];
  assign read_24d[24] = data_0n[24];
  assign read_24d[25] = data_0n[25];
  assign read_24d[26] = data_0n[26];
  assign read_24d[27] = data_0n[27];
  assign read_24d[28] = data_0n[28];
  assign read_24d[29] = data_0n[29];
  assign read_24d[30] = data_0n[30];
  assign read_24d[31] = data_0n[31];
  assign read_24d[32] = data_0n[32];
  assign read_23d[0] = data_0n[0];
  assign read_23d[1] = data_0n[1];
  assign read_23d[2] = data_0n[2];
  assign read_23d[3] = data_0n[3];
  assign read_23d[4] = data_0n[4];
  assign read_23d[5] = data_0n[5];
  assign read_23d[6] = data_0n[6];
  assign read_23d[7] = data_0n[7];
  assign read_23d[8] = data_0n[8];
  assign read_23d[9] = data_0n[9];
  assign read_23d[10] = data_0n[10];
  assign read_23d[11] = data_0n[11];
  assign read_23d[12] = data_0n[12];
  assign read_23d[13] = data_0n[13];
  assign read_23d[14] = data_0n[14];
  assign read_23d[15] = data_0n[15];
  assign read_23d[16] = data_0n[16];
  assign read_23d[17] = data_0n[17];
  assign read_23d[18] = data_0n[18];
  assign read_23d[19] = data_0n[19];
  assign read_23d[20] = data_0n[20];
  assign read_23d[21] = data_0n[21];
  assign read_23d[22] = data_0n[22];
  assign read_23d[23] = data_0n[23];
  assign read_23d[24] = data_0n[24];
  assign read_23d[25] = data_0n[25];
  assign read_23d[26] = data_0n[26];
  assign read_23d[27] = data_0n[27];
  assign read_23d[28] = data_0n[28];
  assign read_23d[29] = data_0n[29];
  assign read_23d[30] = data_0n[30];
  assign read_23d[31] = data_0n[31];
  assign read_23d[32] = data_0n[32];
  assign read_22d[0] = data_0n[0];
  assign read_22d[1] = data_0n[1];
  assign read_22d[2] = data_0n[2];
  assign read_22d[3] = data_0n[3];
  assign read_22d[4] = data_0n[4];
  assign read_22d[5] = data_0n[5];
  assign read_22d[6] = data_0n[6];
  assign read_22d[7] = data_0n[7];
  assign read_22d[8] = data_0n[8];
  assign read_22d[9] = data_0n[9];
  assign read_22d[10] = data_0n[10];
  assign read_22d[11] = data_0n[11];
  assign read_22d[12] = data_0n[12];
  assign read_22d[13] = data_0n[13];
  assign read_22d[14] = data_0n[14];
  assign read_22d[15] = data_0n[15];
  assign read_22d[16] = data_0n[16];
  assign read_22d[17] = data_0n[17];
  assign read_22d[18] = data_0n[18];
  assign read_22d[19] = data_0n[19];
  assign read_22d[20] = data_0n[20];
  assign read_22d[21] = data_0n[21];
  assign read_22d[22] = data_0n[22];
  assign read_22d[23] = data_0n[23];
  assign read_22d[24] = data_0n[24];
  assign read_22d[25] = data_0n[25];
  assign read_22d[26] = data_0n[26];
  assign read_22d[27] = data_0n[27];
  assign read_22d[28] = data_0n[28];
  assign read_22d[29] = data_0n[29];
  assign read_22d[30] = data_0n[30];
  assign read_22d[31] = data_0n[31];
  assign read_22d[32] = data_0n[32];
  assign read_21d[0] = data_0n[0];
  assign read_21d[1] = data_0n[1];
  assign read_21d[2] = data_0n[2];
  assign read_21d[3] = data_0n[3];
  assign read_21d[4] = data_0n[4];
  assign read_21d[5] = data_0n[5];
  assign read_21d[6] = data_0n[6];
  assign read_21d[7] = data_0n[7];
  assign read_21d[8] = data_0n[8];
  assign read_21d[9] = data_0n[9];
  assign read_21d[10] = data_0n[10];
  assign read_21d[11] = data_0n[11];
  assign read_21d[12] = data_0n[12];
  assign read_21d[13] = data_0n[13];
  assign read_21d[14] = data_0n[14];
  assign read_21d[15] = data_0n[15];
  assign read_21d[16] = data_0n[16];
  assign read_21d[17] = data_0n[17];
  assign read_21d[18] = data_0n[18];
  assign read_21d[19] = data_0n[19];
  assign read_21d[20] = data_0n[20];
  assign read_21d[21] = data_0n[21];
  assign read_21d[22] = data_0n[22];
  assign read_21d[23] = data_0n[23];
  assign read_21d[24] = data_0n[24];
  assign read_21d[25] = data_0n[25];
  assign read_21d[26] = data_0n[26];
  assign read_21d[27] = data_0n[27];
  assign read_21d[28] = data_0n[28];
  assign read_21d[29] = data_0n[29];
  assign read_21d[30] = data_0n[30];
  assign read_21d[31] = data_0n[31];
  assign read_21d[32] = data_0n[32];
  assign read_20d[0] = data_0n[0];
  assign read_20d[1] = data_0n[1];
  assign read_20d[2] = data_0n[2];
  assign read_20d[3] = data_0n[3];
  assign read_20d[4] = data_0n[4];
  assign read_20d[5] = data_0n[5];
  assign read_20d[6] = data_0n[6];
  assign read_20d[7] = data_0n[7];
  assign read_20d[8] = data_0n[8];
  assign read_20d[9] = data_0n[9];
  assign read_20d[10] = data_0n[10];
  assign read_20d[11] = data_0n[11];
  assign read_20d[12] = data_0n[12];
  assign read_20d[13] = data_0n[13];
  assign read_20d[14] = data_0n[14];
  assign read_20d[15] = data_0n[15];
  assign read_20d[16] = data_0n[16];
  assign read_20d[17] = data_0n[17];
  assign read_20d[18] = data_0n[18];
  assign read_20d[19] = data_0n[19];
  assign read_20d[20] = data_0n[20];
  assign read_20d[21] = data_0n[21];
  assign read_20d[22] = data_0n[22];
  assign read_20d[23] = data_0n[23];
  assign read_20d[24] = data_0n[24];
  assign read_20d[25] = data_0n[25];
  assign read_20d[26] = data_0n[26];
  assign read_20d[27] = data_0n[27];
  assign read_20d[28] = data_0n[28];
  assign read_20d[29] = data_0n[29];
  assign read_20d[30] = data_0n[30];
  assign read_20d[31] = data_0n[31];
  assign read_20d[32] = data_0n[32];
  assign read_19d[0] = data_0n[0];
  assign read_19d[1] = data_0n[1];
  assign read_19d[2] = data_0n[2];
  assign read_19d[3] = data_0n[3];
  assign read_19d[4] = data_0n[4];
  assign read_19d[5] = data_0n[5];
  assign read_19d[6] = data_0n[6];
  assign read_19d[7] = data_0n[7];
  assign read_19d[8] = data_0n[8];
  assign read_19d[9] = data_0n[9];
  assign read_19d[10] = data_0n[10];
  assign read_19d[11] = data_0n[11];
  assign read_19d[12] = data_0n[12];
  assign read_19d[13] = data_0n[13];
  assign read_19d[14] = data_0n[14];
  assign read_19d[15] = data_0n[15];
  assign read_19d[16] = data_0n[16];
  assign read_19d[17] = data_0n[17];
  assign read_19d[18] = data_0n[18];
  assign read_19d[19] = data_0n[19];
  assign read_19d[20] = data_0n[20];
  assign read_19d[21] = data_0n[21];
  assign read_19d[22] = data_0n[22];
  assign read_19d[23] = data_0n[23];
  assign read_19d[24] = data_0n[24];
  assign read_19d[25] = data_0n[25];
  assign read_19d[26] = data_0n[26];
  assign read_19d[27] = data_0n[27];
  assign read_19d[28] = data_0n[28];
  assign read_19d[29] = data_0n[29];
  assign read_19d[30] = data_0n[30];
  assign read_19d[31] = data_0n[31];
  assign read_19d[32] = data_0n[32];
  assign read_18d[0] = data_0n[0];
  assign read_18d[1] = data_0n[1];
  assign read_18d[2] = data_0n[2];
  assign read_18d[3] = data_0n[3];
  assign read_18d[4] = data_0n[4];
  assign read_18d[5] = data_0n[5];
  assign read_18d[6] = data_0n[6];
  assign read_18d[7] = data_0n[7];
  assign read_18d[8] = data_0n[8];
  assign read_18d[9] = data_0n[9];
  assign read_18d[10] = data_0n[10];
  assign read_18d[11] = data_0n[11];
  assign read_18d[12] = data_0n[12];
  assign read_18d[13] = data_0n[13];
  assign read_18d[14] = data_0n[14];
  assign read_18d[15] = data_0n[15];
  assign read_18d[16] = data_0n[16];
  assign read_18d[17] = data_0n[17];
  assign read_18d[18] = data_0n[18];
  assign read_18d[19] = data_0n[19];
  assign read_18d[20] = data_0n[20];
  assign read_18d[21] = data_0n[21];
  assign read_18d[22] = data_0n[22];
  assign read_18d[23] = data_0n[23];
  assign read_18d[24] = data_0n[24];
  assign read_18d[25] = data_0n[25];
  assign read_18d[26] = data_0n[26];
  assign read_18d[27] = data_0n[27];
  assign read_18d[28] = data_0n[28];
  assign read_18d[29] = data_0n[29];
  assign read_18d[30] = data_0n[30];
  assign read_18d[31] = data_0n[31];
  assign read_18d[32] = data_0n[32];
  assign read_17d[0] = data_0n[0];
  assign read_17d[1] = data_0n[1];
  assign read_17d[2] = data_0n[2];
  assign read_17d[3] = data_0n[3];
  assign read_17d[4] = data_0n[4];
  assign read_17d[5] = data_0n[5];
  assign read_17d[6] = data_0n[6];
  assign read_17d[7] = data_0n[7];
  assign read_17d[8] = data_0n[8];
  assign read_17d[9] = data_0n[9];
  assign read_17d[10] = data_0n[10];
  assign read_17d[11] = data_0n[11];
  assign read_17d[12] = data_0n[12];
  assign read_17d[13] = data_0n[13];
  assign read_17d[14] = data_0n[14];
  assign read_17d[15] = data_0n[15];
  assign read_17d[16] = data_0n[16];
  assign read_17d[17] = data_0n[17];
  assign read_17d[18] = data_0n[18];
  assign read_17d[19] = data_0n[19];
  assign read_17d[20] = data_0n[20];
  assign read_17d[21] = data_0n[21];
  assign read_17d[22] = data_0n[22];
  assign read_17d[23] = data_0n[23];
  assign read_17d[24] = data_0n[24];
  assign read_17d[25] = data_0n[25];
  assign read_17d[26] = data_0n[26];
  assign read_17d[27] = data_0n[27];
  assign read_17d[28] = data_0n[28];
  assign read_17d[29] = data_0n[29];
  assign read_17d[30] = data_0n[30];
  assign read_17d[31] = data_0n[31];
  assign read_17d[32] = data_0n[32];
  assign read_16d[0] = data_0n[0];
  assign read_16d[1] = data_0n[1];
  assign read_16d[2] = data_0n[2];
  assign read_16d[3] = data_0n[3];
  assign read_16d[4] = data_0n[4];
  assign read_16d[5] = data_0n[5];
  assign read_16d[6] = data_0n[6];
  assign read_16d[7] = data_0n[7];
  assign read_16d[8] = data_0n[8];
  assign read_16d[9] = data_0n[9];
  assign read_16d[10] = data_0n[10];
  assign read_16d[11] = data_0n[11];
  assign read_16d[12] = data_0n[12];
  assign read_16d[13] = data_0n[13];
  assign read_16d[14] = data_0n[14];
  assign read_16d[15] = data_0n[15];
  assign read_16d[16] = data_0n[16];
  assign read_16d[17] = data_0n[17];
  assign read_16d[18] = data_0n[18];
  assign read_16d[19] = data_0n[19];
  assign read_16d[20] = data_0n[20];
  assign read_16d[21] = data_0n[21];
  assign read_16d[22] = data_0n[22];
  assign read_16d[23] = data_0n[23];
  assign read_16d[24] = data_0n[24];
  assign read_16d[25] = data_0n[25];
  assign read_16d[26] = data_0n[26];
  assign read_16d[27] = data_0n[27];
  assign read_16d[28] = data_0n[28];
  assign read_16d[29] = data_0n[29];
  assign read_16d[30] = data_0n[30];
  assign read_16d[31] = data_0n[31];
  assign read_16d[32] = data_0n[32];
  assign read_15d[0] = data_0n[0];
  assign read_15d[1] = data_0n[1];
  assign read_15d[2] = data_0n[2];
  assign read_15d[3] = data_0n[3];
  assign read_15d[4] = data_0n[4];
  assign read_15d[5] = data_0n[5];
  assign read_15d[6] = data_0n[6];
  assign read_15d[7] = data_0n[7];
  assign read_15d[8] = data_0n[8];
  assign read_15d[9] = data_0n[9];
  assign read_15d[10] = data_0n[10];
  assign read_15d[11] = data_0n[11];
  assign read_15d[12] = data_0n[12];
  assign read_15d[13] = data_0n[13];
  assign read_15d[14] = data_0n[14];
  assign read_15d[15] = data_0n[15];
  assign read_15d[16] = data_0n[16];
  assign read_15d[17] = data_0n[17];
  assign read_15d[18] = data_0n[18];
  assign read_15d[19] = data_0n[19];
  assign read_15d[20] = data_0n[20];
  assign read_15d[21] = data_0n[21];
  assign read_15d[22] = data_0n[22];
  assign read_15d[23] = data_0n[23];
  assign read_15d[24] = data_0n[24];
  assign read_15d[25] = data_0n[25];
  assign read_15d[26] = data_0n[26];
  assign read_15d[27] = data_0n[27];
  assign read_15d[28] = data_0n[28];
  assign read_15d[29] = data_0n[29];
  assign read_15d[30] = data_0n[30];
  assign read_15d[31] = data_0n[31];
  assign read_15d[32] = data_0n[32];
  assign read_14d[0] = data_0n[0];
  assign read_14d[1] = data_0n[1];
  assign read_14d[2] = data_0n[2];
  assign read_14d[3] = data_0n[3];
  assign read_14d[4] = data_0n[4];
  assign read_14d[5] = data_0n[5];
  assign read_14d[6] = data_0n[6];
  assign read_14d[7] = data_0n[7];
  assign read_14d[8] = data_0n[8];
  assign read_14d[9] = data_0n[9];
  assign read_14d[10] = data_0n[10];
  assign read_14d[11] = data_0n[11];
  assign read_14d[12] = data_0n[12];
  assign read_14d[13] = data_0n[13];
  assign read_14d[14] = data_0n[14];
  assign read_14d[15] = data_0n[15];
  assign read_14d[16] = data_0n[16];
  assign read_14d[17] = data_0n[17];
  assign read_14d[18] = data_0n[18];
  assign read_14d[19] = data_0n[19];
  assign read_14d[20] = data_0n[20];
  assign read_14d[21] = data_0n[21];
  assign read_14d[22] = data_0n[22];
  assign read_14d[23] = data_0n[23];
  assign read_14d[24] = data_0n[24];
  assign read_14d[25] = data_0n[25];
  assign read_14d[26] = data_0n[26];
  assign read_14d[27] = data_0n[27];
  assign read_14d[28] = data_0n[28];
  assign read_14d[29] = data_0n[29];
  assign read_14d[30] = data_0n[30];
  assign read_14d[31] = data_0n[31];
  assign read_14d[32] = data_0n[32];
  assign read_13d[0] = data_0n[0];
  assign read_13d[1] = data_0n[1];
  assign read_13d[2] = data_0n[2];
  assign read_13d[3] = data_0n[3];
  assign read_13d[4] = data_0n[4];
  assign read_13d[5] = data_0n[5];
  assign read_13d[6] = data_0n[6];
  assign read_13d[7] = data_0n[7];
  assign read_13d[8] = data_0n[8];
  assign read_13d[9] = data_0n[9];
  assign read_13d[10] = data_0n[10];
  assign read_13d[11] = data_0n[11];
  assign read_13d[12] = data_0n[12];
  assign read_13d[13] = data_0n[13];
  assign read_13d[14] = data_0n[14];
  assign read_13d[15] = data_0n[15];
  assign read_13d[16] = data_0n[16];
  assign read_13d[17] = data_0n[17];
  assign read_13d[18] = data_0n[18];
  assign read_13d[19] = data_0n[19];
  assign read_13d[20] = data_0n[20];
  assign read_13d[21] = data_0n[21];
  assign read_13d[22] = data_0n[22];
  assign read_13d[23] = data_0n[23];
  assign read_13d[24] = data_0n[24];
  assign read_13d[25] = data_0n[25];
  assign read_13d[26] = data_0n[26];
  assign read_13d[27] = data_0n[27];
  assign read_13d[28] = data_0n[28];
  assign read_13d[29] = data_0n[29];
  assign read_13d[30] = data_0n[30];
  assign read_13d[31] = data_0n[31];
  assign read_13d[32] = data_0n[32];
  assign read_12d[0] = data_0n[0];
  assign read_12d[1] = data_0n[1];
  assign read_12d[2] = data_0n[2];
  assign read_12d[3] = data_0n[3];
  assign read_12d[4] = data_0n[4];
  assign read_12d[5] = data_0n[5];
  assign read_12d[6] = data_0n[6];
  assign read_12d[7] = data_0n[7];
  assign read_12d[8] = data_0n[8];
  assign read_12d[9] = data_0n[9];
  assign read_12d[10] = data_0n[10];
  assign read_12d[11] = data_0n[11];
  assign read_12d[12] = data_0n[12];
  assign read_12d[13] = data_0n[13];
  assign read_12d[14] = data_0n[14];
  assign read_12d[15] = data_0n[15];
  assign read_12d[16] = data_0n[16];
  assign read_12d[17] = data_0n[17];
  assign read_12d[18] = data_0n[18];
  assign read_12d[19] = data_0n[19];
  assign read_12d[20] = data_0n[20];
  assign read_12d[21] = data_0n[21];
  assign read_12d[22] = data_0n[22];
  assign read_12d[23] = data_0n[23];
  assign read_12d[24] = data_0n[24];
  assign read_12d[25] = data_0n[25];
  assign read_12d[26] = data_0n[26];
  assign read_12d[27] = data_0n[27];
  assign read_12d[28] = data_0n[28];
  assign read_12d[29] = data_0n[29];
  assign read_12d[30] = data_0n[30];
  assign read_12d[31] = data_0n[31];
  assign read_12d[32] = data_0n[32];
  assign read_11d[0] = data_0n[0];
  assign read_11d[1] = data_0n[1];
  assign read_11d[2] = data_0n[2];
  assign read_11d[3] = data_0n[3];
  assign read_11d[4] = data_0n[4];
  assign read_11d[5] = data_0n[5];
  assign read_11d[6] = data_0n[6];
  assign read_11d[7] = data_0n[7];
  assign read_11d[8] = data_0n[8];
  assign read_11d[9] = data_0n[9];
  assign read_11d[10] = data_0n[10];
  assign read_11d[11] = data_0n[11];
  assign read_11d[12] = data_0n[12];
  assign read_11d[13] = data_0n[13];
  assign read_11d[14] = data_0n[14];
  assign read_11d[15] = data_0n[15];
  assign read_11d[16] = data_0n[16];
  assign read_11d[17] = data_0n[17];
  assign read_11d[18] = data_0n[18];
  assign read_11d[19] = data_0n[19];
  assign read_11d[20] = data_0n[20];
  assign read_11d[21] = data_0n[21];
  assign read_11d[22] = data_0n[22];
  assign read_11d[23] = data_0n[23];
  assign read_11d[24] = data_0n[24];
  assign read_11d[25] = data_0n[25];
  assign read_11d[26] = data_0n[26];
  assign read_11d[27] = data_0n[27];
  assign read_11d[28] = data_0n[28];
  assign read_11d[29] = data_0n[29];
  assign read_11d[30] = data_0n[30];
  assign read_11d[31] = data_0n[31];
  assign read_11d[32] = data_0n[32];
  assign read_10d[0] = data_0n[0];
  assign read_10d[1] = data_0n[1];
  assign read_10d[2] = data_0n[2];
  assign read_10d[3] = data_0n[3];
  assign read_10d[4] = data_0n[4];
  assign read_10d[5] = data_0n[5];
  assign read_10d[6] = data_0n[6];
  assign read_10d[7] = data_0n[7];
  assign read_10d[8] = data_0n[8];
  assign read_10d[9] = data_0n[9];
  assign read_10d[10] = data_0n[10];
  assign read_10d[11] = data_0n[11];
  assign read_10d[12] = data_0n[12];
  assign read_10d[13] = data_0n[13];
  assign read_10d[14] = data_0n[14];
  assign read_10d[15] = data_0n[15];
  assign read_10d[16] = data_0n[16];
  assign read_10d[17] = data_0n[17];
  assign read_10d[18] = data_0n[18];
  assign read_10d[19] = data_0n[19];
  assign read_10d[20] = data_0n[20];
  assign read_10d[21] = data_0n[21];
  assign read_10d[22] = data_0n[22];
  assign read_10d[23] = data_0n[23];
  assign read_10d[24] = data_0n[24];
  assign read_10d[25] = data_0n[25];
  assign read_10d[26] = data_0n[26];
  assign read_10d[27] = data_0n[27];
  assign read_10d[28] = data_0n[28];
  assign read_10d[29] = data_0n[29];
  assign read_10d[30] = data_0n[30];
  assign read_10d[31] = data_0n[31];
  assign read_10d[32] = data_0n[32];
  assign read_9d[0] = data_0n[0];
  assign read_9d[1] = data_0n[1];
  assign read_9d[2] = data_0n[2];
  assign read_9d[3] = data_0n[3];
  assign read_9d[4] = data_0n[4];
  assign read_9d[5] = data_0n[5];
  assign read_9d[6] = data_0n[6];
  assign read_9d[7] = data_0n[7];
  assign read_9d[8] = data_0n[8];
  assign read_9d[9] = data_0n[9];
  assign read_9d[10] = data_0n[10];
  assign read_9d[11] = data_0n[11];
  assign read_9d[12] = data_0n[12];
  assign read_9d[13] = data_0n[13];
  assign read_9d[14] = data_0n[14];
  assign read_9d[15] = data_0n[15];
  assign read_9d[16] = data_0n[16];
  assign read_9d[17] = data_0n[17];
  assign read_9d[18] = data_0n[18];
  assign read_9d[19] = data_0n[19];
  assign read_9d[20] = data_0n[20];
  assign read_9d[21] = data_0n[21];
  assign read_9d[22] = data_0n[22];
  assign read_9d[23] = data_0n[23];
  assign read_9d[24] = data_0n[24];
  assign read_9d[25] = data_0n[25];
  assign read_9d[26] = data_0n[26];
  assign read_9d[27] = data_0n[27];
  assign read_9d[28] = data_0n[28];
  assign read_9d[29] = data_0n[29];
  assign read_9d[30] = data_0n[30];
  assign read_9d[31] = data_0n[31];
  assign read_9d[32] = data_0n[32];
  assign read_8d[0] = data_0n[0];
  assign read_8d[1] = data_0n[1];
  assign read_8d[2] = data_0n[2];
  assign read_8d[3] = data_0n[3];
  assign read_8d[4] = data_0n[4];
  assign read_8d[5] = data_0n[5];
  assign read_8d[6] = data_0n[6];
  assign read_8d[7] = data_0n[7];
  assign read_8d[8] = data_0n[8];
  assign read_8d[9] = data_0n[9];
  assign read_8d[10] = data_0n[10];
  assign read_8d[11] = data_0n[11];
  assign read_8d[12] = data_0n[12];
  assign read_8d[13] = data_0n[13];
  assign read_8d[14] = data_0n[14];
  assign read_8d[15] = data_0n[15];
  assign read_8d[16] = data_0n[16];
  assign read_8d[17] = data_0n[17];
  assign read_8d[18] = data_0n[18];
  assign read_8d[19] = data_0n[19];
  assign read_8d[20] = data_0n[20];
  assign read_8d[21] = data_0n[21];
  assign read_8d[22] = data_0n[22];
  assign read_8d[23] = data_0n[23];
  assign read_8d[24] = data_0n[24];
  assign read_8d[25] = data_0n[25];
  assign read_8d[26] = data_0n[26];
  assign read_8d[27] = data_0n[27];
  assign read_8d[28] = data_0n[28];
  assign read_8d[29] = data_0n[29];
  assign read_8d[30] = data_0n[30];
  assign read_8d[31] = data_0n[31];
  assign read_8d[32] = data_0n[32];
  assign read_7d[0] = data_0n[0];
  assign read_7d[1] = data_0n[1];
  assign read_7d[2] = data_0n[2];
  assign read_7d[3] = data_0n[3];
  assign read_7d[4] = data_0n[4];
  assign read_7d[5] = data_0n[5];
  assign read_7d[6] = data_0n[6];
  assign read_7d[7] = data_0n[7];
  assign read_7d[8] = data_0n[8];
  assign read_7d[9] = data_0n[9];
  assign read_7d[10] = data_0n[10];
  assign read_7d[11] = data_0n[11];
  assign read_7d[12] = data_0n[12];
  assign read_7d[13] = data_0n[13];
  assign read_7d[14] = data_0n[14];
  assign read_7d[15] = data_0n[15];
  assign read_7d[16] = data_0n[16];
  assign read_7d[17] = data_0n[17];
  assign read_7d[18] = data_0n[18];
  assign read_7d[19] = data_0n[19];
  assign read_7d[20] = data_0n[20];
  assign read_7d[21] = data_0n[21];
  assign read_7d[22] = data_0n[22];
  assign read_7d[23] = data_0n[23];
  assign read_7d[24] = data_0n[24];
  assign read_7d[25] = data_0n[25];
  assign read_7d[26] = data_0n[26];
  assign read_7d[27] = data_0n[27];
  assign read_7d[28] = data_0n[28];
  assign read_7d[29] = data_0n[29];
  assign read_7d[30] = data_0n[30];
  assign read_7d[31] = data_0n[31];
  assign read_7d[32] = data_0n[32];
  assign read_6d[0] = data_0n[0];
  assign read_6d[1] = data_0n[1];
  assign read_6d[2] = data_0n[2];
  assign read_6d[3] = data_0n[3];
  assign read_6d[4] = data_0n[4];
  assign read_6d[5] = data_0n[5];
  assign read_6d[6] = data_0n[6];
  assign read_6d[7] = data_0n[7];
  assign read_6d[8] = data_0n[8];
  assign read_6d[9] = data_0n[9];
  assign read_6d[10] = data_0n[10];
  assign read_6d[11] = data_0n[11];
  assign read_6d[12] = data_0n[12];
  assign read_6d[13] = data_0n[13];
  assign read_6d[14] = data_0n[14];
  assign read_6d[15] = data_0n[15];
  assign read_6d[16] = data_0n[16];
  assign read_6d[17] = data_0n[17];
  assign read_6d[18] = data_0n[18];
  assign read_6d[19] = data_0n[19];
  assign read_6d[20] = data_0n[20];
  assign read_6d[21] = data_0n[21];
  assign read_6d[22] = data_0n[22];
  assign read_6d[23] = data_0n[23];
  assign read_6d[24] = data_0n[24];
  assign read_6d[25] = data_0n[25];
  assign read_6d[26] = data_0n[26];
  assign read_6d[27] = data_0n[27];
  assign read_6d[28] = data_0n[28];
  assign read_6d[29] = data_0n[29];
  assign read_6d[30] = data_0n[30];
  assign read_6d[31] = data_0n[31];
  assign read_6d[32] = data_0n[32];
  assign read_5d[0] = data_0n[0];
  assign read_5d[1] = data_0n[1];
  assign read_5d[2] = data_0n[2];
  assign read_5d[3] = data_0n[3];
  assign read_5d[4] = data_0n[4];
  assign read_5d[5] = data_0n[5];
  assign read_5d[6] = data_0n[6];
  assign read_5d[7] = data_0n[7];
  assign read_5d[8] = data_0n[8];
  assign read_5d[9] = data_0n[9];
  assign read_5d[10] = data_0n[10];
  assign read_5d[11] = data_0n[11];
  assign read_5d[12] = data_0n[12];
  assign read_5d[13] = data_0n[13];
  assign read_5d[14] = data_0n[14];
  assign read_5d[15] = data_0n[15];
  assign read_5d[16] = data_0n[16];
  assign read_5d[17] = data_0n[17];
  assign read_5d[18] = data_0n[18];
  assign read_5d[19] = data_0n[19];
  assign read_5d[20] = data_0n[20];
  assign read_5d[21] = data_0n[21];
  assign read_5d[22] = data_0n[22];
  assign read_5d[23] = data_0n[23];
  assign read_5d[24] = data_0n[24];
  assign read_5d[25] = data_0n[25];
  assign read_5d[26] = data_0n[26];
  assign read_5d[27] = data_0n[27];
  assign read_5d[28] = data_0n[28];
  assign read_5d[29] = data_0n[29];
  assign read_5d[30] = data_0n[30];
  assign read_5d[31] = data_0n[31];
  assign read_5d[32] = data_0n[32];
  assign read_4d[0] = data_0n[0];
  assign read_4d[1] = data_0n[1];
  assign read_4d[2] = data_0n[2];
  assign read_4d[3] = data_0n[3];
  assign read_4d[4] = data_0n[4];
  assign read_4d[5] = data_0n[5];
  assign read_4d[6] = data_0n[6];
  assign read_4d[7] = data_0n[7];
  assign read_4d[8] = data_0n[8];
  assign read_4d[9] = data_0n[9];
  assign read_4d[10] = data_0n[10];
  assign read_4d[11] = data_0n[11];
  assign read_4d[12] = data_0n[12];
  assign read_4d[13] = data_0n[13];
  assign read_4d[14] = data_0n[14];
  assign read_4d[15] = data_0n[15];
  assign read_4d[16] = data_0n[16];
  assign read_4d[17] = data_0n[17];
  assign read_4d[18] = data_0n[18];
  assign read_4d[19] = data_0n[19];
  assign read_4d[20] = data_0n[20];
  assign read_4d[21] = data_0n[21];
  assign read_4d[22] = data_0n[22];
  assign read_4d[23] = data_0n[23];
  assign read_4d[24] = data_0n[24];
  assign read_4d[25] = data_0n[25];
  assign read_4d[26] = data_0n[26];
  assign read_4d[27] = data_0n[27];
  assign read_4d[28] = data_0n[28];
  assign read_4d[29] = data_0n[29];
  assign read_4d[30] = data_0n[30];
  assign read_4d[31] = data_0n[31];
  assign read_4d[32] = data_0n[32];
  assign read_3d[0] = data_0n[0];
  assign read_3d[1] = data_0n[1];
  assign read_3d[2] = data_0n[2];
  assign read_3d[3] = data_0n[3];
  assign read_3d[4] = data_0n[4];
  assign read_3d[5] = data_0n[5];
  assign read_3d[6] = data_0n[6];
  assign read_3d[7] = data_0n[7];
  assign read_3d[8] = data_0n[8];
  assign read_3d[9] = data_0n[9];
  assign read_3d[10] = data_0n[10];
  assign read_3d[11] = data_0n[11];
  assign read_3d[12] = data_0n[12];
  assign read_3d[13] = data_0n[13];
  assign read_3d[14] = data_0n[14];
  assign read_3d[15] = data_0n[15];
  assign read_3d[16] = data_0n[16];
  assign read_3d[17] = data_0n[17];
  assign read_3d[18] = data_0n[18];
  assign read_3d[19] = data_0n[19];
  assign read_3d[20] = data_0n[20];
  assign read_3d[21] = data_0n[21];
  assign read_3d[22] = data_0n[22];
  assign read_3d[23] = data_0n[23];
  assign read_3d[24] = data_0n[24];
  assign read_3d[25] = data_0n[25];
  assign read_3d[26] = data_0n[26];
  assign read_3d[27] = data_0n[27];
  assign read_3d[28] = data_0n[28];
  assign read_3d[29] = data_0n[29];
  assign read_3d[30] = data_0n[30];
  assign read_3d[31] = data_0n[31];
  assign read_3d[32] = data_0n[32];
  assign read_2d[0] = data_0n[0];
  assign read_2d[1] = data_0n[1];
  assign read_2d[2] = data_0n[2];
  assign read_2d[3] = data_0n[3];
  assign read_2d[4] = data_0n[4];
  assign read_2d[5] = data_0n[5];
  assign read_2d[6] = data_0n[6];
  assign read_2d[7] = data_0n[7];
  assign read_2d[8] = data_0n[8];
  assign read_2d[9] = data_0n[9];
  assign read_2d[10] = data_0n[10];
  assign read_2d[11] = data_0n[11];
  assign read_2d[12] = data_0n[12];
  assign read_2d[13] = data_0n[13];
  assign read_2d[14] = data_0n[14];
  assign read_2d[15] = data_0n[15];
  assign read_2d[16] = data_0n[16];
  assign read_2d[17] = data_0n[17];
  assign read_2d[18] = data_0n[18];
  assign read_2d[19] = data_0n[19];
  assign read_2d[20] = data_0n[20];
  assign read_2d[21] = data_0n[21];
  assign read_2d[22] = data_0n[22];
  assign read_2d[23] = data_0n[23];
  assign read_2d[24] = data_0n[24];
  assign read_2d[25] = data_0n[25];
  assign read_2d[26] = data_0n[26];
  assign read_2d[27] = data_0n[27];
  assign read_2d[28] = data_0n[28];
  assign read_2d[29] = data_0n[29];
  assign read_2d[30] = data_0n[30];
  assign read_2d[31] = data_0n[31];
  assign read_2d[32] = data_0n[32];
  assign read_1d[0] = data_0n[0];
  assign read_1d[1] = data_0n[1];
  assign read_1d[2] = data_0n[2];
  assign read_1d[3] = data_0n[3];
  assign read_1d[4] = data_0n[4];
  assign read_1d[5] = data_0n[5];
  assign read_1d[6] = data_0n[6];
  assign read_1d[7] = data_0n[7];
  assign read_1d[8] = data_0n[8];
  assign read_1d[9] = data_0n[9];
  assign read_1d[10] = data_0n[10];
  assign read_1d[11] = data_0n[11];
  assign read_1d[12] = data_0n[12];
  assign read_1d[13] = data_0n[13];
  assign read_1d[14] = data_0n[14];
  assign read_1d[15] = data_0n[15];
  assign read_1d[16] = data_0n[16];
  assign read_1d[17] = data_0n[17];
  assign read_1d[18] = data_0n[18];
  assign read_1d[19] = data_0n[19];
  assign read_1d[20] = data_0n[20];
  assign read_1d[21] = data_0n[21];
  assign read_1d[22] = data_0n[22];
  assign read_1d[23] = data_0n[23];
  assign read_1d[24] = data_0n[24];
  assign read_1d[25] = data_0n[25];
  assign read_1d[26] = data_0n[26];
  assign read_1d[27] = data_0n[27];
  assign read_1d[28] = data_0n[28];
  assign read_1d[29] = data_0n[29];
  assign read_1d[30] = data_0n[30];
  assign read_1d[31] = data_0n[31];
  assign read_1d[32] = data_0n[32];
  assign read_0d[0] = data_0n[0];
  assign read_0d[1] = data_0n[1];
  assign read_0d[2] = data_0n[2];
  assign read_0d[3] = data_0n[3];
  assign read_0d[4] = data_0n[4];
  assign read_0d[5] = data_0n[5];
  assign read_0d[6] = data_0n[6];
  assign read_0d[7] = data_0n[7];
  assign read_0d[8] = data_0n[8];
  assign read_0d[9] = data_0n[9];
  assign read_0d[10] = data_0n[10];
  assign read_0d[11] = data_0n[11];
  assign read_0d[12] = data_0n[12];
  assign read_0d[13] = data_0n[13];
  assign read_0d[14] = data_0n[14];
  assign read_0d[15] = data_0n[15];
  assign read_0d[16] = data_0n[16];
  assign read_0d[17] = data_0n[17];
  assign read_0d[18] = data_0n[18];
  assign read_0d[19] = data_0n[19];
  assign read_0d[20] = data_0n[20];
  assign read_0d[21] = data_0n[21];
  assign read_0d[22] = data_0n[22];
  assign read_0d[23] = data_0n[23];
  assign read_0d[24] = data_0n[24];
  assign read_0d[25] = data_0n[25];
  assign read_0d[26] = data_0n[26];
  assign read_0d[27] = data_0n[27];
  assign read_0d[28] = data_0n[28];
  assign read_0d[29] = data_0n[29];
  assign read_0d[30] = data_0n[30];
  assign read_0d[31] = data_0n[31];
  assign read_0d[32] = data_0n[32];
  LD1 I1088 (write_0d[0], bWriteReq_0n, data_0n[0]);
  LD1 I1089 (write_0d[1], bWriteReq_0n, data_0n[1]);
  LD1 I1090 (write_0d[2], bWriteReq_0n, data_0n[2]);
  LD1 I1091 (write_0d[3], bWriteReq_0n, data_0n[3]);
  LD1 I1092 (write_0d[4], bWriteReq_0n, data_0n[4]);
  LD1 I1093 (write_0d[5], bWriteReq_0n, data_0n[5]);
  LD1 I1094 (write_0d[6], bWriteReq_0n, data_0n[6]);
  LD1 I1095 (write_0d[7], bWriteReq_0n, data_0n[7]);
  LD1 I1096 (write_0d[8], bWriteReq_0n, data_0n[8]);
  LD1 I1097 (write_0d[9], bWriteReq_0n, data_0n[9]);
  LD1 I1098 (write_0d[10], bWriteReq_0n, data_0n[10]);
  LD1 I1099 (write_0d[11], bWriteReq_0n, data_0n[11]);
  LD1 I1100 (write_0d[12], bWriteReq_0n, data_0n[12]);
  LD1 I1101 (write_0d[13], bWriteReq_0n, data_0n[13]);
  LD1 I1102 (write_0d[14], bWriteReq_0n, data_0n[14]);
  LD1 I1103 (write_0d[15], bWriteReq_0n, data_0n[15]);
  LD1 I1104 (write_0d[16], bWriteReq_0n, data_0n[16]);
  LD1 I1105 (write_0d[17], bWriteReq_0n, data_0n[17]);
  LD1 I1106 (write_0d[18], bWriteReq_0n, data_0n[18]);
  LD1 I1107 (write_0d[19], bWriteReq_0n, data_0n[19]);
  LD1 I1108 (write_0d[20], bWriteReq_0n, data_0n[20]);
  LD1 I1109 (write_0d[21], bWriteReq_0n, data_0n[21]);
  LD1 I1110 (write_0d[22], bWriteReq_0n, data_0n[22]);
  LD1 I1111 (write_0d[23], bWriteReq_0n, data_0n[23]);
  LD1 I1112 (write_0d[24], bWriteReq_0n, data_0n[24]);
  LD1 I1113 (write_0d[25], bWriteReq_0n, data_0n[25]);
  LD1 I1114 (write_0d[26], bWriteReq_0n, data_0n[26]);
  LD1 I1115 (write_0d[27], bWriteReq_0n, data_0n[27]);
  LD1 I1116 (write_0d[28], bWriteReq_0n, data_0n[28]);
  LD1 I1117 (write_0d[29], bWriteReq_0n, data_0n[29]);
  LD1 I1118 (write_0d[30], bWriteReq_0n, data_0n[30]);
  LD1 I1119 (write_0d[31], bWriteReq_0n, data_0n[31]);
  LD1 I1120 (write_0d[32], bWriteReq_0n, data_0n[32]);
  IV I1121 (write_0a, nbWriteReq_0n);
  IV I1122 (nbWriteReq_0n, bWriteReq_0n);
  IV I1123 (bWriteReq_0n, nWriteReq_0n);
  IV I1124 (nWriteReq_0n, write_0r);
endmodule

module BrzVariable_33_161_s1305_1_2e_2e1_3b0_2e_2_m4m (
  write_0r, write_0a, write_0d,
  read_0r, read_0a, read_0d,
  read_1r, read_1a, read_1d,
  read_2r, read_2a, read_2d,
  read_3r, read_3a, read_3d,
  read_4r, read_4a, read_4d,
  read_5r, read_5a, read_5d,
  read_6r, read_6a, read_6d,
  read_7r, read_7a, read_7d,
  read_8r, read_8a, read_8d,
  read_9r, read_9a, read_9d,
  read_10r, read_10a, read_10d,
  read_11r, read_11a, read_11d,
  read_12r, read_12a, read_12d,
  read_13r, read_13a, read_13d,
  read_14r, read_14a, read_14d,
  read_15r, read_15a, read_15d,
  read_16r, read_16a, read_16d,
  read_17r, read_17a, read_17d,
  read_18r, read_18a, read_18d,
  read_19r, read_19a, read_19d,
  read_20r, read_20a, read_20d,
  read_21r, read_21a, read_21d,
  read_22r, read_22a, read_22d,
  read_23r, read_23a, read_23d,
  read_24r, read_24a, read_24d,
  read_25r, read_25a, read_25d,
  read_26r, read_26a, read_26d,
  read_27r, read_27a, read_27d,
  read_28r, read_28a, read_28d,
  read_29r, read_29a, read_29d,
  read_30r, read_30a, read_30d,
  read_31r, read_31a, read_31d,
  read_32r, read_32a, read_32d,
  read_33r, read_33a, read_33d,
  read_34r, read_34a, read_34d,
  read_35r, read_35a, read_35d,
  read_36r, read_36a, read_36d,
  read_37r, read_37a, read_37d,
  read_38r, read_38a, read_38d,
  read_39r, read_39a, read_39d,
  read_40r, read_40a, read_40d,
  read_41r, read_41a, read_41d,
  read_42r, read_42a, read_42d,
  read_43r, read_43a, read_43d,
  read_44r, read_44a, read_44d,
  read_45r, read_45a, read_45d,
  read_46r, read_46a, read_46d,
  read_47r, read_47a, read_47d,
  read_48r, read_48a, read_48d,
  read_49r, read_49a, read_49d,
  read_50r, read_50a, read_50d,
  read_51r, read_51a, read_51d,
  read_52r, read_52a, read_52d,
  read_53r, read_53a, read_53d,
  read_54r, read_54a, read_54d,
  read_55r, read_55a, read_55d,
  read_56r, read_56a, read_56d,
  read_57r, read_57a, read_57d,
  read_58r, read_58a, read_58d,
  read_59r, read_59a, read_59d,
  read_60r, read_60a, read_60d,
  read_61r, read_61a, read_61d,
  read_62r, read_62a, read_62d,
  read_63r, read_63a, read_63d,
  read_64r, read_64a, read_64d,
  read_65r, read_65a, read_65d,
  read_66r, read_66a, read_66d,
  read_67r, read_67a, read_67d,
  read_68r, read_68a, read_68d,
  read_69r, read_69a, read_69d,
  read_70r, read_70a, read_70d,
  read_71r, read_71a, read_71d,
  read_72r, read_72a, read_72d,
  read_73r, read_73a, read_73d,
  read_74r, read_74a, read_74d,
  read_75r, read_75a, read_75d,
  read_76r, read_76a, read_76d,
  read_77r, read_77a, read_77d,
  read_78r, read_78a, read_78d,
  read_79r, read_79a, read_79d,
  read_80r, read_80a, read_80d,
  read_81r, read_81a, read_81d,
  read_82r, read_82a, read_82d,
  read_83r, read_83a, read_83d,
  read_84r, read_84a, read_84d,
  read_85r, read_85a, read_85d,
  read_86r, read_86a, read_86d,
  read_87r, read_87a, read_87d,
  read_88r, read_88a, read_88d,
  read_89r, read_89a, read_89d,
  read_90r, read_90a, read_90d,
  read_91r, read_91a, read_91d,
  read_92r, read_92a, read_92d,
  read_93r, read_93a, read_93d,
  read_94r, read_94a, read_94d,
  read_95r, read_95a, read_95d,
  read_96r, read_96a, read_96d,
  read_97r, read_97a, read_97d,
  read_98r, read_98a, read_98d,
  read_99r, read_99a, read_99d,
  read_100r, read_100a, read_100d,
  read_101r, read_101a, read_101d,
  read_102r, read_102a, read_102d,
  read_103r, read_103a, read_103d,
  read_104r, read_104a, read_104d,
  read_105r, read_105a, read_105d,
  read_106r, read_106a, read_106d,
  read_107r, read_107a, read_107d,
  read_108r, read_108a, read_108d,
  read_109r, read_109a, read_109d,
  read_110r, read_110a, read_110d,
  read_111r, read_111a, read_111d,
  read_112r, read_112a, read_112d,
  read_113r, read_113a, read_113d,
  read_114r, read_114a, read_114d,
  read_115r, read_115a, read_115d,
  read_116r, read_116a, read_116d,
  read_117r, read_117a, read_117d,
  read_118r, read_118a, read_118d,
  read_119r, read_119a, read_119d,
  read_120r, read_120a, read_120d,
  read_121r, read_121a, read_121d,
  read_122r, read_122a, read_122d,
  read_123r, read_123a, read_123d,
  read_124r, read_124a, read_124d,
  read_125r, read_125a, read_125d,
  read_126r, read_126a, read_126d,
  read_127r, read_127a, read_127d,
  read_128r, read_128a, read_128d,
  read_129r, read_129a, read_129d,
  read_130r, read_130a, read_130d,
  read_131r, read_131a, read_131d,
  read_132r, read_132a, read_132d,
  read_133r, read_133a, read_133d,
  read_134r, read_134a, read_134d,
  read_135r, read_135a, read_135d,
  read_136r, read_136a, read_136d,
  read_137r, read_137a, read_137d,
  read_138r, read_138a, read_138d,
  read_139r, read_139a, read_139d,
  read_140r, read_140a, read_140d,
  read_141r, read_141a, read_141d,
  read_142r, read_142a, read_142d,
  read_143r, read_143a, read_143d,
  read_144r, read_144a, read_144d,
  read_145r, read_145a, read_145d,
  read_146r, read_146a, read_146d,
  read_147r, read_147a, read_147d,
  read_148r, read_148a, read_148d,
  read_149r, read_149a, read_149d,
  read_150r, read_150a, read_150d,
  read_151r, read_151a, read_151d,
  read_152r, read_152a, read_152d,
  read_153r, read_153a, read_153d,
  read_154r, read_154a, read_154d,
  read_155r, read_155a, read_155d,
  read_156r, read_156a, read_156d,
  read_157r, read_157a, read_157d,
  read_158r, read_158a, read_158d,
  read_159r, read_159a, read_159d,
  read_160r, read_160a, read_160d
);
  input write_0r;
  output write_0a;
  input [32:0] write_0d;
  input read_0r;
  output read_0a;
  output read_0d;
  input read_1r;
  output read_1a;
  output read_1d;
  input read_2r;
  output read_2a;
  output read_2d;
  input read_3r;
  output read_3a;
  output read_3d;
  input read_4r;
  output read_4a;
  output [32:0] read_4d;
  input read_5r;
  output read_5a;
  output [32:0] read_5d;
  input read_6r;
  output read_6a;
  output [32:0] read_6d;
  input read_7r;
  output read_7a;
  output [32:0] read_7d;
  input read_8r;
  output read_8a;
  output [31:0] read_8d;
  input read_9r;
  output read_9a;
  output read_9d;
  input read_10r;
  output read_10a;
  output read_10d;
  input read_11r;
  output read_11a;
  output read_11d;
  input read_12r;
  output read_12a;
  output read_12d;
  input read_13r;
  output read_13a;
  output read_13d;
  input read_14r;
  output read_14a;
  output [32:0] read_14d;
  input read_15r;
  output read_15a;
  output [32:0] read_15d;
  input read_16r;
  output read_16a;
  output [32:0] read_16d;
  input read_17r;
  output read_17a;
  output [32:0] read_17d;
  input read_18r;
  output read_18a;
  output [31:0] read_18d;
  input read_19r;
  output read_19a;
  output read_19d;
  input read_20r;
  output read_20a;
  output read_20d;
  input read_21r;
  output read_21a;
  output read_21d;
  input read_22r;
  output read_22a;
  output read_22d;
  input read_23r;
  output read_23a;
  output read_23d;
  input read_24r;
  output read_24a;
  output [32:0] read_24d;
  input read_25r;
  output read_25a;
  output [32:0] read_25d;
  input read_26r;
  output read_26a;
  output [32:0] read_26d;
  input read_27r;
  output read_27a;
  output [32:0] read_27d;
  input read_28r;
  output read_28a;
  output [31:0] read_28d;
  input read_29r;
  output read_29a;
  output read_29d;
  input read_30r;
  output read_30a;
  output read_30d;
  input read_31r;
  output read_31a;
  output read_31d;
  input read_32r;
  output read_32a;
  output read_32d;
  input read_33r;
  output read_33a;
  output read_33d;
  input read_34r;
  output read_34a;
  output [32:0] read_34d;
  input read_35r;
  output read_35a;
  output [32:0] read_35d;
  input read_36r;
  output read_36a;
  output [32:0] read_36d;
  input read_37r;
  output read_37a;
  output [32:0] read_37d;
  input read_38r;
  output read_38a;
  output [31:0] read_38d;
  input read_39r;
  output read_39a;
  output read_39d;
  input read_40r;
  output read_40a;
  output read_40d;
  input read_41r;
  output read_41a;
  output read_41d;
  input read_42r;
  output read_42a;
  output read_42d;
  input read_43r;
  output read_43a;
  output read_43d;
  input read_44r;
  output read_44a;
  output [32:0] read_44d;
  input read_45r;
  output read_45a;
  output [32:0] read_45d;
  input read_46r;
  output read_46a;
  output [32:0] read_46d;
  input read_47r;
  output read_47a;
  output [32:0] read_47d;
  input read_48r;
  output read_48a;
  output [31:0] read_48d;
  input read_49r;
  output read_49a;
  output read_49d;
  input read_50r;
  output read_50a;
  output read_50d;
  input read_51r;
  output read_51a;
  output read_51d;
  input read_52r;
  output read_52a;
  output read_52d;
  input read_53r;
  output read_53a;
  output read_53d;
  input read_54r;
  output read_54a;
  output [32:0] read_54d;
  input read_55r;
  output read_55a;
  output [32:0] read_55d;
  input read_56r;
  output read_56a;
  output [32:0] read_56d;
  input read_57r;
  output read_57a;
  output [32:0] read_57d;
  input read_58r;
  output read_58a;
  output [31:0] read_58d;
  input read_59r;
  output read_59a;
  output read_59d;
  input read_60r;
  output read_60a;
  output read_60d;
  input read_61r;
  output read_61a;
  output read_61d;
  input read_62r;
  output read_62a;
  output read_62d;
  input read_63r;
  output read_63a;
  output read_63d;
  input read_64r;
  output read_64a;
  output [32:0] read_64d;
  input read_65r;
  output read_65a;
  output [32:0] read_65d;
  input read_66r;
  output read_66a;
  output [32:0] read_66d;
  input read_67r;
  output read_67a;
  output [32:0] read_67d;
  input read_68r;
  output read_68a;
  output [31:0] read_68d;
  input read_69r;
  output read_69a;
  output read_69d;
  input read_70r;
  output read_70a;
  output read_70d;
  input read_71r;
  output read_71a;
  output read_71d;
  input read_72r;
  output read_72a;
  output read_72d;
  input read_73r;
  output read_73a;
  output read_73d;
  input read_74r;
  output read_74a;
  output [32:0] read_74d;
  input read_75r;
  output read_75a;
  output [32:0] read_75d;
  input read_76r;
  output read_76a;
  output [32:0] read_76d;
  input read_77r;
  output read_77a;
  output [32:0] read_77d;
  input read_78r;
  output read_78a;
  output [31:0] read_78d;
  input read_79r;
  output read_79a;
  output read_79d;
  input read_80r;
  output read_80a;
  output read_80d;
  input read_81r;
  output read_81a;
  output read_81d;
  input read_82r;
  output read_82a;
  output read_82d;
  input read_83r;
  output read_83a;
  output read_83d;
  input read_84r;
  output read_84a;
  output [32:0] read_84d;
  input read_85r;
  output read_85a;
  output [32:0] read_85d;
  input read_86r;
  output read_86a;
  output [32:0] read_86d;
  input read_87r;
  output read_87a;
  output [32:0] read_87d;
  input read_88r;
  output read_88a;
  output [31:0] read_88d;
  input read_89r;
  output read_89a;
  output read_89d;
  input read_90r;
  output read_90a;
  output read_90d;
  input read_91r;
  output read_91a;
  output read_91d;
  input read_92r;
  output read_92a;
  output read_92d;
  input read_93r;
  output read_93a;
  output read_93d;
  input read_94r;
  output read_94a;
  output [32:0] read_94d;
  input read_95r;
  output read_95a;
  output [32:0] read_95d;
  input read_96r;
  output read_96a;
  output [32:0] read_96d;
  input read_97r;
  output read_97a;
  output [32:0] read_97d;
  input read_98r;
  output read_98a;
  output [31:0] read_98d;
  input read_99r;
  output read_99a;
  output read_99d;
  input read_100r;
  output read_100a;
  output read_100d;
  input read_101r;
  output read_101a;
  output read_101d;
  input read_102r;
  output read_102a;
  output read_102d;
  input read_103r;
  output read_103a;
  output read_103d;
  input read_104r;
  output read_104a;
  output [32:0] read_104d;
  input read_105r;
  output read_105a;
  output [32:0] read_105d;
  input read_106r;
  output read_106a;
  output [32:0] read_106d;
  input read_107r;
  output read_107a;
  output [32:0] read_107d;
  input read_108r;
  output read_108a;
  output [31:0] read_108d;
  input read_109r;
  output read_109a;
  output read_109d;
  input read_110r;
  output read_110a;
  output read_110d;
  input read_111r;
  output read_111a;
  output read_111d;
  input read_112r;
  output read_112a;
  output read_112d;
  input read_113r;
  output read_113a;
  output read_113d;
  input read_114r;
  output read_114a;
  output [32:0] read_114d;
  input read_115r;
  output read_115a;
  output [32:0] read_115d;
  input read_116r;
  output read_116a;
  output [32:0] read_116d;
  input read_117r;
  output read_117a;
  output [32:0] read_117d;
  input read_118r;
  output read_118a;
  output [31:0] read_118d;
  input read_119r;
  output read_119a;
  output read_119d;
  input read_120r;
  output read_120a;
  output read_120d;
  input read_121r;
  output read_121a;
  output read_121d;
  input read_122r;
  output read_122a;
  output read_122d;
  input read_123r;
  output read_123a;
  output read_123d;
  input read_124r;
  output read_124a;
  output [32:0] read_124d;
  input read_125r;
  output read_125a;
  output [32:0] read_125d;
  input read_126r;
  output read_126a;
  output [32:0] read_126d;
  input read_127r;
  output read_127a;
  output [32:0] read_127d;
  input read_128r;
  output read_128a;
  output [31:0] read_128d;
  input read_129r;
  output read_129a;
  output read_129d;
  input read_130r;
  output read_130a;
  output read_130d;
  input read_131r;
  output read_131a;
  output read_131d;
  input read_132r;
  output read_132a;
  output read_132d;
  input read_133r;
  output read_133a;
  output read_133d;
  input read_134r;
  output read_134a;
  output [32:0] read_134d;
  input read_135r;
  output read_135a;
  output [32:0] read_135d;
  input read_136r;
  output read_136a;
  output [32:0] read_136d;
  input read_137r;
  output read_137a;
  output [32:0] read_137d;
  input read_138r;
  output read_138a;
  output [31:0] read_138d;
  input read_139r;
  output read_139a;
  output read_139d;
  input read_140r;
  output read_140a;
  output read_140d;
  input read_141r;
  output read_141a;
  output read_141d;
  input read_142r;
  output read_142a;
  output read_142d;
  input read_143r;
  output read_143a;
  output read_143d;
  input read_144r;
  output read_144a;
  output [32:0] read_144d;
  input read_145r;
  output read_145a;
  output [32:0] read_145d;
  input read_146r;
  output read_146a;
  output [32:0] read_146d;
  input read_147r;
  output read_147a;
  output [32:0] read_147d;
  input read_148r;
  output read_148a;
  output [31:0] read_148d;
  input read_149r;
  output read_149a;
  output read_149d;
  input read_150r;
  output read_150a;
  output read_150d;
  input read_151r;
  output read_151a;
  output read_151d;
  input read_152r;
  output read_152a;
  output read_152d;
  input read_153r;
  output read_153a;
  output read_153d;
  input read_154r;
  output read_154a;
  output [32:0] read_154d;
  input read_155r;
  output read_155a;
  output [32:0] read_155d;
  input read_156r;
  output read_156a;
  output [32:0] read_156d;
  input read_157r;
  output read_157a;
  output [32:0] read_157d;
  input read_158r;
  output read_158a;
  output [31:0] read_158d;
  input read_159r;
  output read_159a;
  output read_159d;
  input read_160r;
  output read_160a;
  output [31:0] read_160d;
  wire [32:0] data_0n;
  wire nWriteReq_0n;
  wire bWriteReq_0n;
  wire nbWriteReq_0n;
  assign read_0a = read_0r;
  assign read_1a = read_1r;
  assign read_2a = read_2r;
  assign read_3a = read_3r;
  assign read_4a = read_4r;
  assign read_5a = read_5r;
  assign read_6a = read_6r;
  assign read_7a = read_7r;
  assign read_8a = read_8r;
  assign read_9a = read_9r;
  assign read_10a = read_10r;
  assign read_11a = read_11r;
  assign read_12a = read_12r;
  assign read_13a = read_13r;
  assign read_14a = read_14r;
  assign read_15a = read_15r;
  assign read_16a = read_16r;
  assign read_17a = read_17r;
  assign read_18a = read_18r;
  assign read_19a = read_19r;
  assign read_20a = read_20r;
  assign read_21a = read_21r;
  assign read_22a = read_22r;
  assign read_23a = read_23r;
  assign read_24a = read_24r;
  assign read_25a = read_25r;
  assign read_26a = read_26r;
  assign read_27a = read_27r;
  assign read_28a = read_28r;
  assign read_29a = read_29r;
  assign read_30a = read_30r;
  assign read_31a = read_31r;
  assign read_32a = read_32r;
  assign read_33a = read_33r;
  assign read_34a = read_34r;
  assign read_35a = read_35r;
  assign read_36a = read_36r;
  assign read_37a = read_37r;
  assign read_38a = read_38r;
  assign read_39a = read_39r;
  assign read_40a = read_40r;
  assign read_41a = read_41r;
  assign read_42a = read_42r;
  assign read_43a = read_43r;
  assign read_44a = read_44r;
  assign read_45a = read_45r;
  assign read_46a = read_46r;
  assign read_47a = read_47r;
  assign read_48a = read_48r;
  assign read_49a = read_49r;
  assign read_50a = read_50r;
  assign read_51a = read_51r;
  assign read_52a = read_52r;
  assign read_53a = read_53r;
  assign read_54a = read_54r;
  assign read_55a = read_55r;
  assign read_56a = read_56r;
  assign read_57a = read_57r;
  assign read_58a = read_58r;
  assign read_59a = read_59r;
  assign read_60a = read_60r;
  assign read_61a = read_61r;
  assign read_62a = read_62r;
  assign read_63a = read_63r;
  assign read_64a = read_64r;
  assign read_65a = read_65r;
  assign read_66a = read_66r;
  assign read_67a = read_67r;
  assign read_68a = read_68r;
  assign read_69a = read_69r;
  assign read_70a = read_70r;
  assign read_71a = read_71r;
  assign read_72a = read_72r;
  assign read_73a = read_73r;
  assign read_74a = read_74r;
  assign read_75a = read_75r;
  assign read_76a = read_76r;
  assign read_77a = read_77r;
  assign read_78a = read_78r;
  assign read_79a = read_79r;
  assign read_80a = read_80r;
  assign read_81a = read_81r;
  assign read_82a = read_82r;
  assign read_83a = read_83r;
  assign read_84a = read_84r;
  assign read_85a = read_85r;
  assign read_86a = read_86r;
  assign read_87a = read_87r;
  assign read_88a = read_88r;
  assign read_89a = read_89r;
  assign read_90a = read_90r;
  assign read_91a = read_91r;
  assign read_92a = read_92r;
  assign read_93a = read_93r;
  assign read_94a = read_94r;
  assign read_95a = read_95r;
  assign read_96a = read_96r;
  assign read_97a = read_97r;
  assign read_98a = read_98r;
  assign read_99a = read_99r;
  assign read_100a = read_100r;
  assign read_101a = read_101r;
  assign read_102a = read_102r;
  assign read_103a = read_103r;
  assign read_104a = read_104r;
  assign read_105a = read_105r;
  assign read_106a = read_106r;
  assign read_107a = read_107r;
  assign read_108a = read_108r;
  assign read_109a = read_109r;
  assign read_110a = read_110r;
  assign read_111a = read_111r;
  assign read_112a = read_112r;
  assign read_113a = read_113r;
  assign read_114a = read_114r;
  assign read_115a = read_115r;
  assign read_116a = read_116r;
  assign read_117a = read_117r;
  assign read_118a = read_118r;
  assign read_119a = read_119r;
  assign read_120a = read_120r;
  assign read_121a = read_121r;
  assign read_122a = read_122r;
  assign read_123a = read_123r;
  assign read_124a = read_124r;
  assign read_125a = read_125r;
  assign read_126a = read_126r;
  assign read_127a = read_127r;
  assign read_128a = read_128r;
  assign read_129a = read_129r;
  assign read_130a = read_130r;
  assign read_131a = read_131r;
  assign read_132a = read_132r;
  assign read_133a = read_133r;
  assign read_134a = read_134r;
  assign read_135a = read_135r;
  assign read_136a = read_136r;
  assign read_137a = read_137r;
  assign read_138a = read_138r;
  assign read_139a = read_139r;
  assign read_140a = read_140r;
  assign read_141a = read_141r;
  assign read_142a = read_142r;
  assign read_143a = read_143r;
  assign read_144a = read_144r;
  assign read_145a = read_145r;
  assign read_146a = read_146r;
  assign read_147a = read_147r;
  assign read_148a = read_148r;
  assign read_149a = read_149r;
  assign read_150a = read_150r;
  assign read_151a = read_151r;
  assign read_152a = read_152r;
  assign read_153a = read_153r;
  assign read_154a = read_154r;
  assign read_155a = read_155r;
  assign read_156a = read_156r;
  assign read_157a = read_157r;
  assign read_158a = read_158r;
  assign read_159a = read_159r;
  assign read_160a = read_160r;
  assign read_160d[0] = data_0n[1];
  assign read_160d[1] = data_0n[2];
  assign read_160d[2] = data_0n[3];
  assign read_160d[3] = data_0n[4];
  assign read_160d[4] = data_0n[5];
  assign read_160d[5] = data_0n[6];
  assign read_160d[6] = data_0n[7];
  assign read_160d[7] = data_0n[8];
  assign read_160d[8] = data_0n[9];
  assign read_160d[9] = data_0n[10];
  assign read_160d[10] = data_0n[11];
  assign read_160d[11] = data_0n[12];
  assign read_160d[12] = data_0n[13];
  assign read_160d[13] = data_0n[14];
  assign read_160d[14] = data_0n[15];
  assign read_160d[15] = data_0n[16];
  assign read_160d[16] = data_0n[17];
  assign read_160d[17] = data_0n[18];
  assign read_160d[18] = data_0n[19];
  assign read_160d[19] = data_0n[20];
  assign read_160d[20] = data_0n[21];
  assign read_160d[21] = data_0n[22];
  assign read_160d[22] = data_0n[23];
  assign read_160d[23] = data_0n[24];
  assign read_160d[24] = data_0n[25];
  assign read_160d[25] = data_0n[26];
  assign read_160d[26] = data_0n[27];
  assign read_160d[27] = data_0n[28];
  assign read_160d[28] = data_0n[29];
  assign read_160d[29] = data_0n[30];
  assign read_160d[30] = data_0n[31];
  assign read_160d[31] = data_0n[32];
  assign read_159d = data_0n[32];
  assign read_158d[0] = data_0n[1];
  assign read_158d[1] = data_0n[2];
  assign read_158d[2] = data_0n[3];
  assign read_158d[3] = data_0n[4];
  assign read_158d[4] = data_0n[5];
  assign read_158d[5] = data_0n[6];
  assign read_158d[6] = data_0n[7];
  assign read_158d[7] = data_0n[8];
  assign read_158d[8] = data_0n[9];
  assign read_158d[9] = data_0n[10];
  assign read_158d[10] = data_0n[11];
  assign read_158d[11] = data_0n[12];
  assign read_158d[12] = data_0n[13];
  assign read_158d[13] = data_0n[14];
  assign read_158d[14] = data_0n[15];
  assign read_158d[15] = data_0n[16];
  assign read_158d[16] = data_0n[17];
  assign read_158d[17] = data_0n[18];
  assign read_158d[18] = data_0n[19];
  assign read_158d[19] = data_0n[20];
  assign read_158d[20] = data_0n[21];
  assign read_158d[21] = data_0n[22];
  assign read_158d[22] = data_0n[23];
  assign read_158d[23] = data_0n[24];
  assign read_158d[24] = data_0n[25];
  assign read_158d[25] = data_0n[26];
  assign read_158d[26] = data_0n[27];
  assign read_158d[27] = data_0n[28];
  assign read_158d[28] = data_0n[29];
  assign read_158d[29] = data_0n[30];
  assign read_158d[30] = data_0n[31];
  assign read_158d[31] = data_0n[32];
  assign read_157d[0] = data_0n[0];
  assign read_157d[1] = data_0n[1];
  assign read_157d[2] = data_0n[2];
  assign read_157d[3] = data_0n[3];
  assign read_157d[4] = data_0n[4];
  assign read_157d[5] = data_0n[5];
  assign read_157d[6] = data_0n[6];
  assign read_157d[7] = data_0n[7];
  assign read_157d[8] = data_0n[8];
  assign read_157d[9] = data_0n[9];
  assign read_157d[10] = data_0n[10];
  assign read_157d[11] = data_0n[11];
  assign read_157d[12] = data_0n[12];
  assign read_157d[13] = data_0n[13];
  assign read_157d[14] = data_0n[14];
  assign read_157d[15] = data_0n[15];
  assign read_157d[16] = data_0n[16];
  assign read_157d[17] = data_0n[17];
  assign read_157d[18] = data_0n[18];
  assign read_157d[19] = data_0n[19];
  assign read_157d[20] = data_0n[20];
  assign read_157d[21] = data_0n[21];
  assign read_157d[22] = data_0n[22];
  assign read_157d[23] = data_0n[23];
  assign read_157d[24] = data_0n[24];
  assign read_157d[25] = data_0n[25];
  assign read_157d[26] = data_0n[26];
  assign read_157d[27] = data_0n[27];
  assign read_157d[28] = data_0n[28];
  assign read_157d[29] = data_0n[29];
  assign read_157d[30] = data_0n[30];
  assign read_157d[31] = data_0n[31];
  assign read_157d[32] = data_0n[32];
  assign read_156d[0] = data_0n[0];
  assign read_156d[1] = data_0n[1];
  assign read_156d[2] = data_0n[2];
  assign read_156d[3] = data_0n[3];
  assign read_156d[4] = data_0n[4];
  assign read_156d[5] = data_0n[5];
  assign read_156d[6] = data_0n[6];
  assign read_156d[7] = data_0n[7];
  assign read_156d[8] = data_0n[8];
  assign read_156d[9] = data_0n[9];
  assign read_156d[10] = data_0n[10];
  assign read_156d[11] = data_0n[11];
  assign read_156d[12] = data_0n[12];
  assign read_156d[13] = data_0n[13];
  assign read_156d[14] = data_0n[14];
  assign read_156d[15] = data_0n[15];
  assign read_156d[16] = data_0n[16];
  assign read_156d[17] = data_0n[17];
  assign read_156d[18] = data_0n[18];
  assign read_156d[19] = data_0n[19];
  assign read_156d[20] = data_0n[20];
  assign read_156d[21] = data_0n[21];
  assign read_156d[22] = data_0n[22];
  assign read_156d[23] = data_0n[23];
  assign read_156d[24] = data_0n[24];
  assign read_156d[25] = data_0n[25];
  assign read_156d[26] = data_0n[26];
  assign read_156d[27] = data_0n[27];
  assign read_156d[28] = data_0n[28];
  assign read_156d[29] = data_0n[29];
  assign read_156d[30] = data_0n[30];
  assign read_156d[31] = data_0n[31];
  assign read_156d[32] = data_0n[32];
  assign read_155d[0] = data_0n[0];
  assign read_155d[1] = data_0n[1];
  assign read_155d[2] = data_0n[2];
  assign read_155d[3] = data_0n[3];
  assign read_155d[4] = data_0n[4];
  assign read_155d[5] = data_0n[5];
  assign read_155d[6] = data_0n[6];
  assign read_155d[7] = data_0n[7];
  assign read_155d[8] = data_0n[8];
  assign read_155d[9] = data_0n[9];
  assign read_155d[10] = data_0n[10];
  assign read_155d[11] = data_0n[11];
  assign read_155d[12] = data_0n[12];
  assign read_155d[13] = data_0n[13];
  assign read_155d[14] = data_0n[14];
  assign read_155d[15] = data_0n[15];
  assign read_155d[16] = data_0n[16];
  assign read_155d[17] = data_0n[17];
  assign read_155d[18] = data_0n[18];
  assign read_155d[19] = data_0n[19];
  assign read_155d[20] = data_0n[20];
  assign read_155d[21] = data_0n[21];
  assign read_155d[22] = data_0n[22];
  assign read_155d[23] = data_0n[23];
  assign read_155d[24] = data_0n[24];
  assign read_155d[25] = data_0n[25];
  assign read_155d[26] = data_0n[26];
  assign read_155d[27] = data_0n[27];
  assign read_155d[28] = data_0n[28];
  assign read_155d[29] = data_0n[29];
  assign read_155d[30] = data_0n[30];
  assign read_155d[31] = data_0n[31];
  assign read_155d[32] = data_0n[32];
  assign read_154d[0] = data_0n[0];
  assign read_154d[1] = data_0n[1];
  assign read_154d[2] = data_0n[2];
  assign read_154d[3] = data_0n[3];
  assign read_154d[4] = data_0n[4];
  assign read_154d[5] = data_0n[5];
  assign read_154d[6] = data_0n[6];
  assign read_154d[7] = data_0n[7];
  assign read_154d[8] = data_0n[8];
  assign read_154d[9] = data_0n[9];
  assign read_154d[10] = data_0n[10];
  assign read_154d[11] = data_0n[11];
  assign read_154d[12] = data_0n[12];
  assign read_154d[13] = data_0n[13];
  assign read_154d[14] = data_0n[14];
  assign read_154d[15] = data_0n[15];
  assign read_154d[16] = data_0n[16];
  assign read_154d[17] = data_0n[17];
  assign read_154d[18] = data_0n[18];
  assign read_154d[19] = data_0n[19];
  assign read_154d[20] = data_0n[20];
  assign read_154d[21] = data_0n[21];
  assign read_154d[22] = data_0n[22];
  assign read_154d[23] = data_0n[23];
  assign read_154d[24] = data_0n[24];
  assign read_154d[25] = data_0n[25];
  assign read_154d[26] = data_0n[26];
  assign read_154d[27] = data_0n[27];
  assign read_154d[28] = data_0n[28];
  assign read_154d[29] = data_0n[29];
  assign read_154d[30] = data_0n[30];
  assign read_154d[31] = data_0n[31];
  assign read_154d[32] = data_0n[32];
  assign read_153d = data_0n[0];
  assign read_152d = data_0n[1];
  assign read_151d = data_0n[0];
  assign read_150d = data_0n[1];
  assign read_149d = data_0n[32];
  assign read_148d[0] = data_0n[1];
  assign read_148d[1] = data_0n[2];
  assign read_148d[2] = data_0n[3];
  assign read_148d[3] = data_0n[4];
  assign read_148d[4] = data_0n[5];
  assign read_148d[5] = data_0n[6];
  assign read_148d[6] = data_0n[7];
  assign read_148d[7] = data_0n[8];
  assign read_148d[8] = data_0n[9];
  assign read_148d[9] = data_0n[10];
  assign read_148d[10] = data_0n[11];
  assign read_148d[11] = data_0n[12];
  assign read_148d[12] = data_0n[13];
  assign read_148d[13] = data_0n[14];
  assign read_148d[14] = data_0n[15];
  assign read_148d[15] = data_0n[16];
  assign read_148d[16] = data_0n[17];
  assign read_148d[17] = data_0n[18];
  assign read_148d[18] = data_0n[19];
  assign read_148d[19] = data_0n[20];
  assign read_148d[20] = data_0n[21];
  assign read_148d[21] = data_0n[22];
  assign read_148d[22] = data_0n[23];
  assign read_148d[23] = data_0n[24];
  assign read_148d[24] = data_0n[25];
  assign read_148d[25] = data_0n[26];
  assign read_148d[26] = data_0n[27];
  assign read_148d[27] = data_0n[28];
  assign read_148d[28] = data_0n[29];
  assign read_148d[29] = data_0n[30];
  assign read_148d[30] = data_0n[31];
  assign read_148d[31] = data_0n[32];
  assign read_147d[0] = data_0n[0];
  assign read_147d[1] = data_0n[1];
  assign read_147d[2] = data_0n[2];
  assign read_147d[3] = data_0n[3];
  assign read_147d[4] = data_0n[4];
  assign read_147d[5] = data_0n[5];
  assign read_147d[6] = data_0n[6];
  assign read_147d[7] = data_0n[7];
  assign read_147d[8] = data_0n[8];
  assign read_147d[9] = data_0n[9];
  assign read_147d[10] = data_0n[10];
  assign read_147d[11] = data_0n[11];
  assign read_147d[12] = data_0n[12];
  assign read_147d[13] = data_0n[13];
  assign read_147d[14] = data_0n[14];
  assign read_147d[15] = data_0n[15];
  assign read_147d[16] = data_0n[16];
  assign read_147d[17] = data_0n[17];
  assign read_147d[18] = data_0n[18];
  assign read_147d[19] = data_0n[19];
  assign read_147d[20] = data_0n[20];
  assign read_147d[21] = data_0n[21];
  assign read_147d[22] = data_0n[22];
  assign read_147d[23] = data_0n[23];
  assign read_147d[24] = data_0n[24];
  assign read_147d[25] = data_0n[25];
  assign read_147d[26] = data_0n[26];
  assign read_147d[27] = data_0n[27];
  assign read_147d[28] = data_0n[28];
  assign read_147d[29] = data_0n[29];
  assign read_147d[30] = data_0n[30];
  assign read_147d[31] = data_0n[31];
  assign read_147d[32] = data_0n[32];
  assign read_146d[0] = data_0n[0];
  assign read_146d[1] = data_0n[1];
  assign read_146d[2] = data_0n[2];
  assign read_146d[3] = data_0n[3];
  assign read_146d[4] = data_0n[4];
  assign read_146d[5] = data_0n[5];
  assign read_146d[6] = data_0n[6];
  assign read_146d[7] = data_0n[7];
  assign read_146d[8] = data_0n[8];
  assign read_146d[9] = data_0n[9];
  assign read_146d[10] = data_0n[10];
  assign read_146d[11] = data_0n[11];
  assign read_146d[12] = data_0n[12];
  assign read_146d[13] = data_0n[13];
  assign read_146d[14] = data_0n[14];
  assign read_146d[15] = data_0n[15];
  assign read_146d[16] = data_0n[16];
  assign read_146d[17] = data_0n[17];
  assign read_146d[18] = data_0n[18];
  assign read_146d[19] = data_0n[19];
  assign read_146d[20] = data_0n[20];
  assign read_146d[21] = data_0n[21];
  assign read_146d[22] = data_0n[22];
  assign read_146d[23] = data_0n[23];
  assign read_146d[24] = data_0n[24];
  assign read_146d[25] = data_0n[25];
  assign read_146d[26] = data_0n[26];
  assign read_146d[27] = data_0n[27];
  assign read_146d[28] = data_0n[28];
  assign read_146d[29] = data_0n[29];
  assign read_146d[30] = data_0n[30];
  assign read_146d[31] = data_0n[31];
  assign read_146d[32] = data_0n[32];
  assign read_145d[0] = data_0n[0];
  assign read_145d[1] = data_0n[1];
  assign read_145d[2] = data_0n[2];
  assign read_145d[3] = data_0n[3];
  assign read_145d[4] = data_0n[4];
  assign read_145d[5] = data_0n[5];
  assign read_145d[6] = data_0n[6];
  assign read_145d[7] = data_0n[7];
  assign read_145d[8] = data_0n[8];
  assign read_145d[9] = data_0n[9];
  assign read_145d[10] = data_0n[10];
  assign read_145d[11] = data_0n[11];
  assign read_145d[12] = data_0n[12];
  assign read_145d[13] = data_0n[13];
  assign read_145d[14] = data_0n[14];
  assign read_145d[15] = data_0n[15];
  assign read_145d[16] = data_0n[16];
  assign read_145d[17] = data_0n[17];
  assign read_145d[18] = data_0n[18];
  assign read_145d[19] = data_0n[19];
  assign read_145d[20] = data_0n[20];
  assign read_145d[21] = data_0n[21];
  assign read_145d[22] = data_0n[22];
  assign read_145d[23] = data_0n[23];
  assign read_145d[24] = data_0n[24];
  assign read_145d[25] = data_0n[25];
  assign read_145d[26] = data_0n[26];
  assign read_145d[27] = data_0n[27];
  assign read_145d[28] = data_0n[28];
  assign read_145d[29] = data_0n[29];
  assign read_145d[30] = data_0n[30];
  assign read_145d[31] = data_0n[31];
  assign read_145d[32] = data_0n[32];
  assign read_144d[0] = data_0n[0];
  assign read_144d[1] = data_0n[1];
  assign read_144d[2] = data_0n[2];
  assign read_144d[3] = data_0n[3];
  assign read_144d[4] = data_0n[4];
  assign read_144d[5] = data_0n[5];
  assign read_144d[6] = data_0n[6];
  assign read_144d[7] = data_0n[7];
  assign read_144d[8] = data_0n[8];
  assign read_144d[9] = data_0n[9];
  assign read_144d[10] = data_0n[10];
  assign read_144d[11] = data_0n[11];
  assign read_144d[12] = data_0n[12];
  assign read_144d[13] = data_0n[13];
  assign read_144d[14] = data_0n[14];
  assign read_144d[15] = data_0n[15];
  assign read_144d[16] = data_0n[16];
  assign read_144d[17] = data_0n[17];
  assign read_144d[18] = data_0n[18];
  assign read_144d[19] = data_0n[19];
  assign read_144d[20] = data_0n[20];
  assign read_144d[21] = data_0n[21];
  assign read_144d[22] = data_0n[22];
  assign read_144d[23] = data_0n[23];
  assign read_144d[24] = data_0n[24];
  assign read_144d[25] = data_0n[25];
  assign read_144d[26] = data_0n[26];
  assign read_144d[27] = data_0n[27];
  assign read_144d[28] = data_0n[28];
  assign read_144d[29] = data_0n[29];
  assign read_144d[30] = data_0n[30];
  assign read_144d[31] = data_0n[31];
  assign read_144d[32] = data_0n[32];
  assign read_143d = data_0n[0];
  assign read_142d = data_0n[1];
  assign read_141d = data_0n[0];
  assign read_140d = data_0n[1];
  assign read_139d = data_0n[32];
  assign read_138d[0] = data_0n[1];
  assign read_138d[1] = data_0n[2];
  assign read_138d[2] = data_0n[3];
  assign read_138d[3] = data_0n[4];
  assign read_138d[4] = data_0n[5];
  assign read_138d[5] = data_0n[6];
  assign read_138d[6] = data_0n[7];
  assign read_138d[7] = data_0n[8];
  assign read_138d[8] = data_0n[9];
  assign read_138d[9] = data_0n[10];
  assign read_138d[10] = data_0n[11];
  assign read_138d[11] = data_0n[12];
  assign read_138d[12] = data_0n[13];
  assign read_138d[13] = data_0n[14];
  assign read_138d[14] = data_0n[15];
  assign read_138d[15] = data_0n[16];
  assign read_138d[16] = data_0n[17];
  assign read_138d[17] = data_0n[18];
  assign read_138d[18] = data_0n[19];
  assign read_138d[19] = data_0n[20];
  assign read_138d[20] = data_0n[21];
  assign read_138d[21] = data_0n[22];
  assign read_138d[22] = data_0n[23];
  assign read_138d[23] = data_0n[24];
  assign read_138d[24] = data_0n[25];
  assign read_138d[25] = data_0n[26];
  assign read_138d[26] = data_0n[27];
  assign read_138d[27] = data_0n[28];
  assign read_138d[28] = data_0n[29];
  assign read_138d[29] = data_0n[30];
  assign read_138d[30] = data_0n[31];
  assign read_138d[31] = data_0n[32];
  assign read_137d[0] = data_0n[0];
  assign read_137d[1] = data_0n[1];
  assign read_137d[2] = data_0n[2];
  assign read_137d[3] = data_0n[3];
  assign read_137d[4] = data_0n[4];
  assign read_137d[5] = data_0n[5];
  assign read_137d[6] = data_0n[6];
  assign read_137d[7] = data_0n[7];
  assign read_137d[8] = data_0n[8];
  assign read_137d[9] = data_0n[9];
  assign read_137d[10] = data_0n[10];
  assign read_137d[11] = data_0n[11];
  assign read_137d[12] = data_0n[12];
  assign read_137d[13] = data_0n[13];
  assign read_137d[14] = data_0n[14];
  assign read_137d[15] = data_0n[15];
  assign read_137d[16] = data_0n[16];
  assign read_137d[17] = data_0n[17];
  assign read_137d[18] = data_0n[18];
  assign read_137d[19] = data_0n[19];
  assign read_137d[20] = data_0n[20];
  assign read_137d[21] = data_0n[21];
  assign read_137d[22] = data_0n[22];
  assign read_137d[23] = data_0n[23];
  assign read_137d[24] = data_0n[24];
  assign read_137d[25] = data_0n[25];
  assign read_137d[26] = data_0n[26];
  assign read_137d[27] = data_0n[27];
  assign read_137d[28] = data_0n[28];
  assign read_137d[29] = data_0n[29];
  assign read_137d[30] = data_0n[30];
  assign read_137d[31] = data_0n[31];
  assign read_137d[32] = data_0n[32];
  assign read_136d[0] = data_0n[0];
  assign read_136d[1] = data_0n[1];
  assign read_136d[2] = data_0n[2];
  assign read_136d[3] = data_0n[3];
  assign read_136d[4] = data_0n[4];
  assign read_136d[5] = data_0n[5];
  assign read_136d[6] = data_0n[6];
  assign read_136d[7] = data_0n[7];
  assign read_136d[8] = data_0n[8];
  assign read_136d[9] = data_0n[9];
  assign read_136d[10] = data_0n[10];
  assign read_136d[11] = data_0n[11];
  assign read_136d[12] = data_0n[12];
  assign read_136d[13] = data_0n[13];
  assign read_136d[14] = data_0n[14];
  assign read_136d[15] = data_0n[15];
  assign read_136d[16] = data_0n[16];
  assign read_136d[17] = data_0n[17];
  assign read_136d[18] = data_0n[18];
  assign read_136d[19] = data_0n[19];
  assign read_136d[20] = data_0n[20];
  assign read_136d[21] = data_0n[21];
  assign read_136d[22] = data_0n[22];
  assign read_136d[23] = data_0n[23];
  assign read_136d[24] = data_0n[24];
  assign read_136d[25] = data_0n[25];
  assign read_136d[26] = data_0n[26];
  assign read_136d[27] = data_0n[27];
  assign read_136d[28] = data_0n[28];
  assign read_136d[29] = data_0n[29];
  assign read_136d[30] = data_0n[30];
  assign read_136d[31] = data_0n[31];
  assign read_136d[32] = data_0n[32];
  assign read_135d[0] = data_0n[0];
  assign read_135d[1] = data_0n[1];
  assign read_135d[2] = data_0n[2];
  assign read_135d[3] = data_0n[3];
  assign read_135d[4] = data_0n[4];
  assign read_135d[5] = data_0n[5];
  assign read_135d[6] = data_0n[6];
  assign read_135d[7] = data_0n[7];
  assign read_135d[8] = data_0n[8];
  assign read_135d[9] = data_0n[9];
  assign read_135d[10] = data_0n[10];
  assign read_135d[11] = data_0n[11];
  assign read_135d[12] = data_0n[12];
  assign read_135d[13] = data_0n[13];
  assign read_135d[14] = data_0n[14];
  assign read_135d[15] = data_0n[15];
  assign read_135d[16] = data_0n[16];
  assign read_135d[17] = data_0n[17];
  assign read_135d[18] = data_0n[18];
  assign read_135d[19] = data_0n[19];
  assign read_135d[20] = data_0n[20];
  assign read_135d[21] = data_0n[21];
  assign read_135d[22] = data_0n[22];
  assign read_135d[23] = data_0n[23];
  assign read_135d[24] = data_0n[24];
  assign read_135d[25] = data_0n[25];
  assign read_135d[26] = data_0n[26];
  assign read_135d[27] = data_0n[27];
  assign read_135d[28] = data_0n[28];
  assign read_135d[29] = data_0n[29];
  assign read_135d[30] = data_0n[30];
  assign read_135d[31] = data_0n[31];
  assign read_135d[32] = data_0n[32];
  assign read_134d[0] = data_0n[0];
  assign read_134d[1] = data_0n[1];
  assign read_134d[2] = data_0n[2];
  assign read_134d[3] = data_0n[3];
  assign read_134d[4] = data_0n[4];
  assign read_134d[5] = data_0n[5];
  assign read_134d[6] = data_0n[6];
  assign read_134d[7] = data_0n[7];
  assign read_134d[8] = data_0n[8];
  assign read_134d[9] = data_0n[9];
  assign read_134d[10] = data_0n[10];
  assign read_134d[11] = data_0n[11];
  assign read_134d[12] = data_0n[12];
  assign read_134d[13] = data_0n[13];
  assign read_134d[14] = data_0n[14];
  assign read_134d[15] = data_0n[15];
  assign read_134d[16] = data_0n[16];
  assign read_134d[17] = data_0n[17];
  assign read_134d[18] = data_0n[18];
  assign read_134d[19] = data_0n[19];
  assign read_134d[20] = data_0n[20];
  assign read_134d[21] = data_0n[21];
  assign read_134d[22] = data_0n[22];
  assign read_134d[23] = data_0n[23];
  assign read_134d[24] = data_0n[24];
  assign read_134d[25] = data_0n[25];
  assign read_134d[26] = data_0n[26];
  assign read_134d[27] = data_0n[27];
  assign read_134d[28] = data_0n[28];
  assign read_134d[29] = data_0n[29];
  assign read_134d[30] = data_0n[30];
  assign read_134d[31] = data_0n[31];
  assign read_134d[32] = data_0n[32];
  assign read_133d = data_0n[0];
  assign read_132d = data_0n[1];
  assign read_131d = data_0n[0];
  assign read_130d = data_0n[1];
  assign read_129d = data_0n[32];
  assign read_128d[0] = data_0n[1];
  assign read_128d[1] = data_0n[2];
  assign read_128d[2] = data_0n[3];
  assign read_128d[3] = data_0n[4];
  assign read_128d[4] = data_0n[5];
  assign read_128d[5] = data_0n[6];
  assign read_128d[6] = data_0n[7];
  assign read_128d[7] = data_0n[8];
  assign read_128d[8] = data_0n[9];
  assign read_128d[9] = data_0n[10];
  assign read_128d[10] = data_0n[11];
  assign read_128d[11] = data_0n[12];
  assign read_128d[12] = data_0n[13];
  assign read_128d[13] = data_0n[14];
  assign read_128d[14] = data_0n[15];
  assign read_128d[15] = data_0n[16];
  assign read_128d[16] = data_0n[17];
  assign read_128d[17] = data_0n[18];
  assign read_128d[18] = data_0n[19];
  assign read_128d[19] = data_0n[20];
  assign read_128d[20] = data_0n[21];
  assign read_128d[21] = data_0n[22];
  assign read_128d[22] = data_0n[23];
  assign read_128d[23] = data_0n[24];
  assign read_128d[24] = data_0n[25];
  assign read_128d[25] = data_0n[26];
  assign read_128d[26] = data_0n[27];
  assign read_128d[27] = data_0n[28];
  assign read_128d[28] = data_0n[29];
  assign read_128d[29] = data_0n[30];
  assign read_128d[30] = data_0n[31];
  assign read_128d[31] = data_0n[32];
  assign read_127d[0] = data_0n[0];
  assign read_127d[1] = data_0n[1];
  assign read_127d[2] = data_0n[2];
  assign read_127d[3] = data_0n[3];
  assign read_127d[4] = data_0n[4];
  assign read_127d[5] = data_0n[5];
  assign read_127d[6] = data_0n[6];
  assign read_127d[7] = data_0n[7];
  assign read_127d[8] = data_0n[8];
  assign read_127d[9] = data_0n[9];
  assign read_127d[10] = data_0n[10];
  assign read_127d[11] = data_0n[11];
  assign read_127d[12] = data_0n[12];
  assign read_127d[13] = data_0n[13];
  assign read_127d[14] = data_0n[14];
  assign read_127d[15] = data_0n[15];
  assign read_127d[16] = data_0n[16];
  assign read_127d[17] = data_0n[17];
  assign read_127d[18] = data_0n[18];
  assign read_127d[19] = data_0n[19];
  assign read_127d[20] = data_0n[20];
  assign read_127d[21] = data_0n[21];
  assign read_127d[22] = data_0n[22];
  assign read_127d[23] = data_0n[23];
  assign read_127d[24] = data_0n[24];
  assign read_127d[25] = data_0n[25];
  assign read_127d[26] = data_0n[26];
  assign read_127d[27] = data_0n[27];
  assign read_127d[28] = data_0n[28];
  assign read_127d[29] = data_0n[29];
  assign read_127d[30] = data_0n[30];
  assign read_127d[31] = data_0n[31];
  assign read_127d[32] = data_0n[32];
  assign read_126d[0] = data_0n[0];
  assign read_126d[1] = data_0n[1];
  assign read_126d[2] = data_0n[2];
  assign read_126d[3] = data_0n[3];
  assign read_126d[4] = data_0n[4];
  assign read_126d[5] = data_0n[5];
  assign read_126d[6] = data_0n[6];
  assign read_126d[7] = data_0n[7];
  assign read_126d[8] = data_0n[8];
  assign read_126d[9] = data_0n[9];
  assign read_126d[10] = data_0n[10];
  assign read_126d[11] = data_0n[11];
  assign read_126d[12] = data_0n[12];
  assign read_126d[13] = data_0n[13];
  assign read_126d[14] = data_0n[14];
  assign read_126d[15] = data_0n[15];
  assign read_126d[16] = data_0n[16];
  assign read_126d[17] = data_0n[17];
  assign read_126d[18] = data_0n[18];
  assign read_126d[19] = data_0n[19];
  assign read_126d[20] = data_0n[20];
  assign read_126d[21] = data_0n[21];
  assign read_126d[22] = data_0n[22];
  assign read_126d[23] = data_0n[23];
  assign read_126d[24] = data_0n[24];
  assign read_126d[25] = data_0n[25];
  assign read_126d[26] = data_0n[26];
  assign read_126d[27] = data_0n[27];
  assign read_126d[28] = data_0n[28];
  assign read_126d[29] = data_0n[29];
  assign read_126d[30] = data_0n[30];
  assign read_126d[31] = data_0n[31];
  assign read_126d[32] = data_0n[32];
  assign read_125d[0] = data_0n[0];
  assign read_125d[1] = data_0n[1];
  assign read_125d[2] = data_0n[2];
  assign read_125d[3] = data_0n[3];
  assign read_125d[4] = data_0n[4];
  assign read_125d[5] = data_0n[5];
  assign read_125d[6] = data_0n[6];
  assign read_125d[7] = data_0n[7];
  assign read_125d[8] = data_0n[8];
  assign read_125d[9] = data_0n[9];
  assign read_125d[10] = data_0n[10];
  assign read_125d[11] = data_0n[11];
  assign read_125d[12] = data_0n[12];
  assign read_125d[13] = data_0n[13];
  assign read_125d[14] = data_0n[14];
  assign read_125d[15] = data_0n[15];
  assign read_125d[16] = data_0n[16];
  assign read_125d[17] = data_0n[17];
  assign read_125d[18] = data_0n[18];
  assign read_125d[19] = data_0n[19];
  assign read_125d[20] = data_0n[20];
  assign read_125d[21] = data_0n[21];
  assign read_125d[22] = data_0n[22];
  assign read_125d[23] = data_0n[23];
  assign read_125d[24] = data_0n[24];
  assign read_125d[25] = data_0n[25];
  assign read_125d[26] = data_0n[26];
  assign read_125d[27] = data_0n[27];
  assign read_125d[28] = data_0n[28];
  assign read_125d[29] = data_0n[29];
  assign read_125d[30] = data_0n[30];
  assign read_125d[31] = data_0n[31];
  assign read_125d[32] = data_0n[32];
  assign read_124d[0] = data_0n[0];
  assign read_124d[1] = data_0n[1];
  assign read_124d[2] = data_0n[2];
  assign read_124d[3] = data_0n[3];
  assign read_124d[4] = data_0n[4];
  assign read_124d[5] = data_0n[5];
  assign read_124d[6] = data_0n[6];
  assign read_124d[7] = data_0n[7];
  assign read_124d[8] = data_0n[8];
  assign read_124d[9] = data_0n[9];
  assign read_124d[10] = data_0n[10];
  assign read_124d[11] = data_0n[11];
  assign read_124d[12] = data_0n[12];
  assign read_124d[13] = data_0n[13];
  assign read_124d[14] = data_0n[14];
  assign read_124d[15] = data_0n[15];
  assign read_124d[16] = data_0n[16];
  assign read_124d[17] = data_0n[17];
  assign read_124d[18] = data_0n[18];
  assign read_124d[19] = data_0n[19];
  assign read_124d[20] = data_0n[20];
  assign read_124d[21] = data_0n[21];
  assign read_124d[22] = data_0n[22];
  assign read_124d[23] = data_0n[23];
  assign read_124d[24] = data_0n[24];
  assign read_124d[25] = data_0n[25];
  assign read_124d[26] = data_0n[26];
  assign read_124d[27] = data_0n[27];
  assign read_124d[28] = data_0n[28];
  assign read_124d[29] = data_0n[29];
  assign read_124d[30] = data_0n[30];
  assign read_124d[31] = data_0n[31];
  assign read_124d[32] = data_0n[32];
  assign read_123d = data_0n[0];
  assign read_122d = data_0n[1];
  assign read_121d = data_0n[0];
  assign read_120d = data_0n[1];
  assign read_119d = data_0n[32];
  assign read_118d[0] = data_0n[1];
  assign read_118d[1] = data_0n[2];
  assign read_118d[2] = data_0n[3];
  assign read_118d[3] = data_0n[4];
  assign read_118d[4] = data_0n[5];
  assign read_118d[5] = data_0n[6];
  assign read_118d[6] = data_0n[7];
  assign read_118d[7] = data_0n[8];
  assign read_118d[8] = data_0n[9];
  assign read_118d[9] = data_0n[10];
  assign read_118d[10] = data_0n[11];
  assign read_118d[11] = data_0n[12];
  assign read_118d[12] = data_0n[13];
  assign read_118d[13] = data_0n[14];
  assign read_118d[14] = data_0n[15];
  assign read_118d[15] = data_0n[16];
  assign read_118d[16] = data_0n[17];
  assign read_118d[17] = data_0n[18];
  assign read_118d[18] = data_0n[19];
  assign read_118d[19] = data_0n[20];
  assign read_118d[20] = data_0n[21];
  assign read_118d[21] = data_0n[22];
  assign read_118d[22] = data_0n[23];
  assign read_118d[23] = data_0n[24];
  assign read_118d[24] = data_0n[25];
  assign read_118d[25] = data_0n[26];
  assign read_118d[26] = data_0n[27];
  assign read_118d[27] = data_0n[28];
  assign read_118d[28] = data_0n[29];
  assign read_118d[29] = data_0n[30];
  assign read_118d[30] = data_0n[31];
  assign read_118d[31] = data_0n[32];
  assign read_117d[0] = data_0n[0];
  assign read_117d[1] = data_0n[1];
  assign read_117d[2] = data_0n[2];
  assign read_117d[3] = data_0n[3];
  assign read_117d[4] = data_0n[4];
  assign read_117d[5] = data_0n[5];
  assign read_117d[6] = data_0n[6];
  assign read_117d[7] = data_0n[7];
  assign read_117d[8] = data_0n[8];
  assign read_117d[9] = data_0n[9];
  assign read_117d[10] = data_0n[10];
  assign read_117d[11] = data_0n[11];
  assign read_117d[12] = data_0n[12];
  assign read_117d[13] = data_0n[13];
  assign read_117d[14] = data_0n[14];
  assign read_117d[15] = data_0n[15];
  assign read_117d[16] = data_0n[16];
  assign read_117d[17] = data_0n[17];
  assign read_117d[18] = data_0n[18];
  assign read_117d[19] = data_0n[19];
  assign read_117d[20] = data_0n[20];
  assign read_117d[21] = data_0n[21];
  assign read_117d[22] = data_0n[22];
  assign read_117d[23] = data_0n[23];
  assign read_117d[24] = data_0n[24];
  assign read_117d[25] = data_0n[25];
  assign read_117d[26] = data_0n[26];
  assign read_117d[27] = data_0n[27];
  assign read_117d[28] = data_0n[28];
  assign read_117d[29] = data_0n[29];
  assign read_117d[30] = data_0n[30];
  assign read_117d[31] = data_0n[31];
  assign read_117d[32] = data_0n[32];
  assign read_116d[0] = data_0n[0];
  assign read_116d[1] = data_0n[1];
  assign read_116d[2] = data_0n[2];
  assign read_116d[3] = data_0n[3];
  assign read_116d[4] = data_0n[4];
  assign read_116d[5] = data_0n[5];
  assign read_116d[6] = data_0n[6];
  assign read_116d[7] = data_0n[7];
  assign read_116d[8] = data_0n[8];
  assign read_116d[9] = data_0n[9];
  assign read_116d[10] = data_0n[10];
  assign read_116d[11] = data_0n[11];
  assign read_116d[12] = data_0n[12];
  assign read_116d[13] = data_0n[13];
  assign read_116d[14] = data_0n[14];
  assign read_116d[15] = data_0n[15];
  assign read_116d[16] = data_0n[16];
  assign read_116d[17] = data_0n[17];
  assign read_116d[18] = data_0n[18];
  assign read_116d[19] = data_0n[19];
  assign read_116d[20] = data_0n[20];
  assign read_116d[21] = data_0n[21];
  assign read_116d[22] = data_0n[22];
  assign read_116d[23] = data_0n[23];
  assign read_116d[24] = data_0n[24];
  assign read_116d[25] = data_0n[25];
  assign read_116d[26] = data_0n[26];
  assign read_116d[27] = data_0n[27];
  assign read_116d[28] = data_0n[28];
  assign read_116d[29] = data_0n[29];
  assign read_116d[30] = data_0n[30];
  assign read_116d[31] = data_0n[31];
  assign read_116d[32] = data_0n[32];
  assign read_115d[0] = data_0n[0];
  assign read_115d[1] = data_0n[1];
  assign read_115d[2] = data_0n[2];
  assign read_115d[3] = data_0n[3];
  assign read_115d[4] = data_0n[4];
  assign read_115d[5] = data_0n[5];
  assign read_115d[6] = data_0n[6];
  assign read_115d[7] = data_0n[7];
  assign read_115d[8] = data_0n[8];
  assign read_115d[9] = data_0n[9];
  assign read_115d[10] = data_0n[10];
  assign read_115d[11] = data_0n[11];
  assign read_115d[12] = data_0n[12];
  assign read_115d[13] = data_0n[13];
  assign read_115d[14] = data_0n[14];
  assign read_115d[15] = data_0n[15];
  assign read_115d[16] = data_0n[16];
  assign read_115d[17] = data_0n[17];
  assign read_115d[18] = data_0n[18];
  assign read_115d[19] = data_0n[19];
  assign read_115d[20] = data_0n[20];
  assign read_115d[21] = data_0n[21];
  assign read_115d[22] = data_0n[22];
  assign read_115d[23] = data_0n[23];
  assign read_115d[24] = data_0n[24];
  assign read_115d[25] = data_0n[25];
  assign read_115d[26] = data_0n[26];
  assign read_115d[27] = data_0n[27];
  assign read_115d[28] = data_0n[28];
  assign read_115d[29] = data_0n[29];
  assign read_115d[30] = data_0n[30];
  assign read_115d[31] = data_0n[31];
  assign read_115d[32] = data_0n[32];
  assign read_114d[0] = data_0n[0];
  assign read_114d[1] = data_0n[1];
  assign read_114d[2] = data_0n[2];
  assign read_114d[3] = data_0n[3];
  assign read_114d[4] = data_0n[4];
  assign read_114d[5] = data_0n[5];
  assign read_114d[6] = data_0n[6];
  assign read_114d[7] = data_0n[7];
  assign read_114d[8] = data_0n[8];
  assign read_114d[9] = data_0n[9];
  assign read_114d[10] = data_0n[10];
  assign read_114d[11] = data_0n[11];
  assign read_114d[12] = data_0n[12];
  assign read_114d[13] = data_0n[13];
  assign read_114d[14] = data_0n[14];
  assign read_114d[15] = data_0n[15];
  assign read_114d[16] = data_0n[16];
  assign read_114d[17] = data_0n[17];
  assign read_114d[18] = data_0n[18];
  assign read_114d[19] = data_0n[19];
  assign read_114d[20] = data_0n[20];
  assign read_114d[21] = data_0n[21];
  assign read_114d[22] = data_0n[22];
  assign read_114d[23] = data_0n[23];
  assign read_114d[24] = data_0n[24];
  assign read_114d[25] = data_0n[25];
  assign read_114d[26] = data_0n[26];
  assign read_114d[27] = data_0n[27];
  assign read_114d[28] = data_0n[28];
  assign read_114d[29] = data_0n[29];
  assign read_114d[30] = data_0n[30];
  assign read_114d[31] = data_0n[31];
  assign read_114d[32] = data_0n[32];
  assign read_113d = data_0n[0];
  assign read_112d = data_0n[1];
  assign read_111d = data_0n[0];
  assign read_110d = data_0n[1];
  assign read_109d = data_0n[32];
  assign read_108d[0] = data_0n[1];
  assign read_108d[1] = data_0n[2];
  assign read_108d[2] = data_0n[3];
  assign read_108d[3] = data_0n[4];
  assign read_108d[4] = data_0n[5];
  assign read_108d[5] = data_0n[6];
  assign read_108d[6] = data_0n[7];
  assign read_108d[7] = data_0n[8];
  assign read_108d[8] = data_0n[9];
  assign read_108d[9] = data_0n[10];
  assign read_108d[10] = data_0n[11];
  assign read_108d[11] = data_0n[12];
  assign read_108d[12] = data_0n[13];
  assign read_108d[13] = data_0n[14];
  assign read_108d[14] = data_0n[15];
  assign read_108d[15] = data_0n[16];
  assign read_108d[16] = data_0n[17];
  assign read_108d[17] = data_0n[18];
  assign read_108d[18] = data_0n[19];
  assign read_108d[19] = data_0n[20];
  assign read_108d[20] = data_0n[21];
  assign read_108d[21] = data_0n[22];
  assign read_108d[22] = data_0n[23];
  assign read_108d[23] = data_0n[24];
  assign read_108d[24] = data_0n[25];
  assign read_108d[25] = data_0n[26];
  assign read_108d[26] = data_0n[27];
  assign read_108d[27] = data_0n[28];
  assign read_108d[28] = data_0n[29];
  assign read_108d[29] = data_0n[30];
  assign read_108d[30] = data_0n[31];
  assign read_108d[31] = data_0n[32];
  assign read_107d[0] = data_0n[0];
  assign read_107d[1] = data_0n[1];
  assign read_107d[2] = data_0n[2];
  assign read_107d[3] = data_0n[3];
  assign read_107d[4] = data_0n[4];
  assign read_107d[5] = data_0n[5];
  assign read_107d[6] = data_0n[6];
  assign read_107d[7] = data_0n[7];
  assign read_107d[8] = data_0n[8];
  assign read_107d[9] = data_0n[9];
  assign read_107d[10] = data_0n[10];
  assign read_107d[11] = data_0n[11];
  assign read_107d[12] = data_0n[12];
  assign read_107d[13] = data_0n[13];
  assign read_107d[14] = data_0n[14];
  assign read_107d[15] = data_0n[15];
  assign read_107d[16] = data_0n[16];
  assign read_107d[17] = data_0n[17];
  assign read_107d[18] = data_0n[18];
  assign read_107d[19] = data_0n[19];
  assign read_107d[20] = data_0n[20];
  assign read_107d[21] = data_0n[21];
  assign read_107d[22] = data_0n[22];
  assign read_107d[23] = data_0n[23];
  assign read_107d[24] = data_0n[24];
  assign read_107d[25] = data_0n[25];
  assign read_107d[26] = data_0n[26];
  assign read_107d[27] = data_0n[27];
  assign read_107d[28] = data_0n[28];
  assign read_107d[29] = data_0n[29];
  assign read_107d[30] = data_0n[30];
  assign read_107d[31] = data_0n[31];
  assign read_107d[32] = data_0n[32];
  assign read_106d[0] = data_0n[0];
  assign read_106d[1] = data_0n[1];
  assign read_106d[2] = data_0n[2];
  assign read_106d[3] = data_0n[3];
  assign read_106d[4] = data_0n[4];
  assign read_106d[5] = data_0n[5];
  assign read_106d[6] = data_0n[6];
  assign read_106d[7] = data_0n[7];
  assign read_106d[8] = data_0n[8];
  assign read_106d[9] = data_0n[9];
  assign read_106d[10] = data_0n[10];
  assign read_106d[11] = data_0n[11];
  assign read_106d[12] = data_0n[12];
  assign read_106d[13] = data_0n[13];
  assign read_106d[14] = data_0n[14];
  assign read_106d[15] = data_0n[15];
  assign read_106d[16] = data_0n[16];
  assign read_106d[17] = data_0n[17];
  assign read_106d[18] = data_0n[18];
  assign read_106d[19] = data_0n[19];
  assign read_106d[20] = data_0n[20];
  assign read_106d[21] = data_0n[21];
  assign read_106d[22] = data_0n[22];
  assign read_106d[23] = data_0n[23];
  assign read_106d[24] = data_0n[24];
  assign read_106d[25] = data_0n[25];
  assign read_106d[26] = data_0n[26];
  assign read_106d[27] = data_0n[27];
  assign read_106d[28] = data_0n[28];
  assign read_106d[29] = data_0n[29];
  assign read_106d[30] = data_0n[30];
  assign read_106d[31] = data_0n[31];
  assign read_106d[32] = data_0n[32];
  assign read_105d[0] = data_0n[0];
  assign read_105d[1] = data_0n[1];
  assign read_105d[2] = data_0n[2];
  assign read_105d[3] = data_0n[3];
  assign read_105d[4] = data_0n[4];
  assign read_105d[5] = data_0n[5];
  assign read_105d[6] = data_0n[6];
  assign read_105d[7] = data_0n[7];
  assign read_105d[8] = data_0n[8];
  assign read_105d[9] = data_0n[9];
  assign read_105d[10] = data_0n[10];
  assign read_105d[11] = data_0n[11];
  assign read_105d[12] = data_0n[12];
  assign read_105d[13] = data_0n[13];
  assign read_105d[14] = data_0n[14];
  assign read_105d[15] = data_0n[15];
  assign read_105d[16] = data_0n[16];
  assign read_105d[17] = data_0n[17];
  assign read_105d[18] = data_0n[18];
  assign read_105d[19] = data_0n[19];
  assign read_105d[20] = data_0n[20];
  assign read_105d[21] = data_0n[21];
  assign read_105d[22] = data_0n[22];
  assign read_105d[23] = data_0n[23];
  assign read_105d[24] = data_0n[24];
  assign read_105d[25] = data_0n[25];
  assign read_105d[26] = data_0n[26];
  assign read_105d[27] = data_0n[27];
  assign read_105d[28] = data_0n[28];
  assign read_105d[29] = data_0n[29];
  assign read_105d[30] = data_0n[30];
  assign read_105d[31] = data_0n[31];
  assign read_105d[32] = data_0n[32];
  assign read_104d[0] = data_0n[0];
  assign read_104d[1] = data_0n[1];
  assign read_104d[2] = data_0n[2];
  assign read_104d[3] = data_0n[3];
  assign read_104d[4] = data_0n[4];
  assign read_104d[5] = data_0n[5];
  assign read_104d[6] = data_0n[6];
  assign read_104d[7] = data_0n[7];
  assign read_104d[8] = data_0n[8];
  assign read_104d[9] = data_0n[9];
  assign read_104d[10] = data_0n[10];
  assign read_104d[11] = data_0n[11];
  assign read_104d[12] = data_0n[12];
  assign read_104d[13] = data_0n[13];
  assign read_104d[14] = data_0n[14];
  assign read_104d[15] = data_0n[15];
  assign read_104d[16] = data_0n[16];
  assign read_104d[17] = data_0n[17];
  assign read_104d[18] = data_0n[18];
  assign read_104d[19] = data_0n[19];
  assign read_104d[20] = data_0n[20];
  assign read_104d[21] = data_0n[21];
  assign read_104d[22] = data_0n[22];
  assign read_104d[23] = data_0n[23];
  assign read_104d[24] = data_0n[24];
  assign read_104d[25] = data_0n[25];
  assign read_104d[26] = data_0n[26];
  assign read_104d[27] = data_0n[27];
  assign read_104d[28] = data_0n[28];
  assign read_104d[29] = data_0n[29];
  assign read_104d[30] = data_0n[30];
  assign read_104d[31] = data_0n[31];
  assign read_104d[32] = data_0n[32];
  assign read_103d = data_0n[0];
  assign read_102d = data_0n[1];
  assign read_101d = data_0n[0];
  assign read_100d = data_0n[1];
  assign read_99d = data_0n[32];
  assign read_98d[0] = data_0n[1];
  assign read_98d[1] = data_0n[2];
  assign read_98d[2] = data_0n[3];
  assign read_98d[3] = data_0n[4];
  assign read_98d[4] = data_0n[5];
  assign read_98d[5] = data_0n[6];
  assign read_98d[6] = data_0n[7];
  assign read_98d[7] = data_0n[8];
  assign read_98d[8] = data_0n[9];
  assign read_98d[9] = data_0n[10];
  assign read_98d[10] = data_0n[11];
  assign read_98d[11] = data_0n[12];
  assign read_98d[12] = data_0n[13];
  assign read_98d[13] = data_0n[14];
  assign read_98d[14] = data_0n[15];
  assign read_98d[15] = data_0n[16];
  assign read_98d[16] = data_0n[17];
  assign read_98d[17] = data_0n[18];
  assign read_98d[18] = data_0n[19];
  assign read_98d[19] = data_0n[20];
  assign read_98d[20] = data_0n[21];
  assign read_98d[21] = data_0n[22];
  assign read_98d[22] = data_0n[23];
  assign read_98d[23] = data_0n[24];
  assign read_98d[24] = data_0n[25];
  assign read_98d[25] = data_0n[26];
  assign read_98d[26] = data_0n[27];
  assign read_98d[27] = data_0n[28];
  assign read_98d[28] = data_0n[29];
  assign read_98d[29] = data_0n[30];
  assign read_98d[30] = data_0n[31];
  assign read_98d[31] = data_0n[32];
  assign read_97d[0] = data_0n[0];
  assign read_97d[1] = data_0n[1];
  assign read_97d[2] = data_0n[2];
  assign read_97d[3] = data_0n[3];
  assign read_97d[4] = data_0n[4];
  assign read_97d[5] = data_0n[5];
  assign read_97d[6] = data_0n[6];
  assign read_97d[7] = data_0n[7];
  assign read_97d[8] = data_0n[8];
  assign read_97d[9] = data_0n[9];
  assign read_97d[10] = data_0n[10];
  assign read_97d[11] = data_0n[11];
  assign read_97d[12] = data_0n[12];
  assign read_97d[13] = data_0n[13];
  assign read_97d[14] = data_0n[14];
  assign read_97d[15] = data_0n[15];
  assign read_97d[16] = data_0n[16];
  assign read_97d[17] = data_0n[17];
  assign read_97d[18] = data_0n[18];
  assign read_97d[19] = data_0n[19];
  assign read_97d[20] = data_0n[20];
  assign read_97d[21] = data_0n[21];
  assign read_97d[22] = data_0n[22];
  assign read_97d[23] = data_0n[23];
  assign read_97d[24] = data_0n[24];
  assign read_97d[25] = data_0n[25];
  assign read_97d[26] = data_0n[26];
  assign read_97d[27] = data_0n[27];
  assign read_97d[28] = data_0n[28];
  assign read_97d[29] = data_0n[29];
  assign read_97d[30] = data_0n[30];
  assign read_97d[31] = data_0n[31];
  assign read_97d[32] = data_0n[32];
  assign read_96d[0] = data_0n[0];
  assign read_96d[1] = data_0n[1];
  assign read_96d[2] = data_0n[2];
  assign read_96d[3] = data_0n[3];
  assign read_96d[4] = data_0n[4];
  assign read_96d[5] = data_0n[5];
  assign read_96d[6] = data_0n[6];
  assign read_96d[7] = data_0n[7];
  assign read_96d[8] = data_0n[8];
  assign read_96d[9] = data_0n[9];
  assign read_96d[10] = data_0n[10];
  assign read_96d[11] = data_0n[11];
  assign read_96d[12] = data_0n[12];
  assign read_96d[13] = data_0n[13];
  assign read_96d[14] = data_0n[14];
  assign read_96d[15] = data_0n[15];
  assign read_96d[16] = data_0n[16];
  assign read_96d[17] = data_0n[17];
  assign read_96d[18] = data_0n[18];
  assign read_96d[19] = data_0n[19];
  assign read_96d[20] = data_0n[20];
  assign read_96d[21] = data_0n[21];
  assign read_96d[22] = data_0n[22];
  assign read_96d[23] = data_0n[23];
  assign read_96d[24] = data_0n[24];
  assign read_96d[25] = data_0n[25];
  assign read_96d[26] = data_0n[26];
  assign read_96d[27] = data_0n[27];
  assign read_96d[28] = data_0n[28];
  assign read_96d[29] = data_0n[29];
  assign read_96d[30] = data_0n[30];
  assign read_96d[31] = data_0n[31];
  assign read_96d[32] = data_0n[32];
  assign read_95d[0] = data_0n[0];
  assign read_95d[1] = data_0n[1];
  assign read_95d[2] = data_0n[2];
  assign read_95d[3] = data_0n[3];
  assign read_95d[4] = data_0n[4];
  assign read_95d[5] = data_0n[5];
  assign read_95d[6] = data_0n[6];
  assign read_95d[7] = data_0n[7];
  assign read_95d[8] = data_0n[8];
  assign read_95d[9] = data_0n[9];
  assign read_95d[10] = data_0n[10];
  assign read_95d[11] = data_0n[11];
  assign read_95d[12] = data_0n[12];
  assign read_95d[13] = data_0n[13];
  assign read_95d[14] = data_0n[14];
  assign read_95d[15] = data_0n[15];
  assign read_95d[16] = data_0n[16];
  assign read_95d[17] = data_0n[17];
  assign read_95d[18] = data_0n[18];
  assign read_95d[19] = data_0n[19];
  assign read_95d[20] = data_0n[20];
  assign read_95d[21] = data_0n[21];
  assign read_95d[22] = data_0n[22];
  assign read_95d[23] = data_0n[23];
  assign read_95d[24] = data_0n[24];
  assign read_95d[25] = data_0n[25];
  assign read_95d[26] = data_0n[26];
  assign read_95d[27] = data_0n[27];
  assign read_95d[28] = data_0n[28];
  assign read_95d[29] = data_0n[29];
  assign read_95d[30] = data_0n[30];
  assign read_95d[31] = data_0n[31];
  assign read_95d[32] = data_0n[32];
  assign read_94d[0] = data_0n[0];
  assign read_94d[1] = data_0n[1];
  assign read_94d[2] = data_0n[2];
  assign read_94d[3] = data_0n[3];
  assign read_94d[4] = data_0n[4];
  assign read_94d[5] = data_0n[5];
  assign read_94d[6] = data_0n[6];
  assign read_94d[7] = data_0n[7];
  assign read_94d[8] = data_0n[8];
  assign read_94d[9] = data_0n[9];
  assign read_94d[10] = data_0n[10];
  assign read_94d[11] = data_0n[11];
  assign read_94d[12] = data_0n[12];
  assign read_94d[13] = data_0n[13];
  assign read_94d[14] = data_0n[14];
  assign read_94d[15] = data_0n[15];
  assign read_94d[16] = data_0n[16];
  assign read_94d[17] = data_0n[17];
  assign read_94d[18] = data_0n[18];
  assign read_94d[19] = data_0n[19];
  assign read_94d[20] = data_0n[20];
  assign read_94d[21] = data_0n[21];
  assign read_94d[22] = data_0n[22];
  assign read_94d[23] = data_0n[23];
  assign read_94d[24] = data_0n[24];
  assign read_94d[25] = data_0n[25];
  assign read_94d[26] = data_0n[26];
  assign read_94d[27] = data_0n[27];
  assign read_94d[28] = data_0n[28];
  assign read_94d[29] = data_0n[29];
  assign read_94d[30] = data_0n[30];
  assign read_94d[31] = data_0n[31];
  assign read_94d[32] = data_0n[32];
  assign read_93d = data_0n[0];
  assign read_92d = data_0n[1];
  assign read_91d = data_0n[0];
  assign read_90d = data_0n[1];
  assign read_89d = data_0n[32];
  assign read_88d[0] = data_0n[1];
  assign read_88d[1] = data_0n[2];
  assign read_88d[2] = data_0n[3];
  assign read_88d[3] = data_0n[4];
  assign read_88d[4] = data_0n[5];
  assign read_88d[5] = data_0n[6];
  assign read_88d[6] = data_0n[7];
  assign read_88d[7] = data_0n[8];
  assign read_88d[8] = data_0n[9];
  assign read_88d[9] = data_0n[10];
  assign read_88d[10] = data_0n[11];
  assign read_88d[11] = data_0n[12];
  assign read_88d[12] = data_0n[13];
  assign read_88d[13] = data_0n[14];
  assign read_88d[14] = data_0n[15];
  assign read_88d[15] = data_0n[16];
  assign read_88d[16] = data_0n[17];
  assign read_88d[17] = data_0n[18];
  assign read_88d[18] = data_0n[19];
  assign read_88d[19] = data_0n[20];
  assign read_88d[20] = data_0n[21];
  assign read_88d[21] = data_0n[22];
  assign read_88d[22] = data_0n[23];
  assign read_88d[23] = data_0n[24];
  assign read_88d[24] = data_0n[25];
  assign read_88d[25] = data_0n[26];
  assign read_88d[26] = data_0n[27];
  assign read_88d[27] = data_0n[28];
  assign read_88d[28] = data_0n[29];
  assign read_88d[29] = data_0n[30];
  assign read_88d[30] = data_0n[31];
  assign read_88d[31] = data_0n[32];
  assign read_87d[0] = data_0n[0];
  assign read_87d[1] = data_0n[1];
  assign read_87d[2] = data_0n[2];
  assign read_87d[3] = data_0n[3];
  assign read_87d[4] = data_0n[4];
  assign read_87d[5] = data_0n[5];
  assign read_87d[6] = data_0n[6];
  assign read_87d[7] = data_0n[7];
  assign read_87d[8] = data_0n[8];
  assign read_87d[9] = data_0n[9];
  assign read_87d[10] = data_0n[10];
  assign read_87d[11] = data_0n[11];
  assign read_87d[12] = data_0n[12];
  assign read_87d[13] = data_0n[13];
  assign read_87d[14] = data_0n[14];
  assign read_87d[15] = data_0n[15];
  assign read_87d[16] = data_0n[16];
  assign read_87d[17] = data_0n[17];
  assign read_87d[18] = data_0n[18];
  assign read_87d[19] = data_0n[19];
  assign read_87d[20] = data_0n[20];
  assign read_87d[21] = data_0n[21];
  assign read_87d[22] = data_0n[22];
  assign read_87d[23] = data_0n[23];
  assign read_87d[24] = data_0n[24];
  assign read_87d[25] = data_0n[25];
  assign read_87d[26] = data_0n[26];
  assign read_87d[27] = data_0n[27];
  assign read_87d[28] = data_0n[28];
  assign read_87d[29] = data_0n[29];
  assign read_87d[30] = data_0n[30];
  assign read_87d[31] = data_0n[31];
  assign read_87d[32] = data_0n[32];
  assign read_86d[0] = data_0n[0];
  assign read_86d[1] = data_0n[1];
  assign read_86d[2] = data_0n[2];
  assign read_86d[3] = data_0n[3];
  assign read_86d[4] = data_0n[4];
  assign read_86d[5] = data_0n[5];
  assign read_86d[6] = data_0n[6];
  assign read_86d[7] = data_0n[7];
  assign read_86d[8] = data_0n[8];
  assign read_86d[9] = data_0n[9];
  assign read_86d[10] = data_0n[10];
  assign read_86d[11] = data_0n[11];
  assign read_86d[12] = data_0n[12];
  assign read_86d[13] = data_0n[13];
  assign read_86d[14] = data_0n[14];
  assign read_86d[15] = data_0n[15];
  assign read_86d[16] = data_0n[16];
  assign read_86d[17] = data_0n[17];
  assign read_86d[18] = data_0n[18];
  assign read_86d[19] = data_0n[19];
  assign read_86d[20] = data_0n[20];
  assign read_86d[21] = data_0n[21];
  assign read_86d[22] = data_0n[22];
  assign read_86d[23] = data_0n[23];
  assign read_86d[24] = data_0n[24];
  assign read_86d[25] = data_0n[25];
  assign read_86d[26] = data_0n[26];
  assign read_86d[27] = data_0n[27];
  assign read_86d[28] = data_0n[28];
  assign read_86d[29] = data_0n[29];
  assign read_86d[30] = data_0n[30];
  assign read_86d[31] = data_0n[31];
  assign read_86d[32] = data_0n[32];
  assign read_85d[0] = data_0n[0];
  assign read_85d[1] = data_0n[1];
  assign read_85d[2] = data_0n[2];
  assign read_85d[3] = data_0n[3];
  assign read_85d[4] = data_0n[4];
  assign read_85d[5] = data_0n[5];
  assign read_85d[6] = data_0n[6];
  assign read_85d[7] = data_0n[7];
  assign read_85d[8] = data_0n[8];
  assign read_85d[9] = data_0n[9];
  assign read_85d[10] = data_0n[10];
  assign read_85d[11] = data_0n[11];
  assign read_85d[12] = data_0n[12];
  assign read_85d[13] = data_0n[13];
  assign read_85d[14] = data_0n[14];
  assign read_85d[15] = data_0n[15];
  assign read_85d[16] = data_0n[16];
  assign read_85d[17] = data_0n[17];
  assign read_85d[18] = data_0n[18];
  assign read_85d[19] = data_0n[19];
  assign read_85d[20] = data_0n[20];
  assign read_85d[21] = data_0n[21];
  assign read_85d[22] = data_0n[22];
  assign read_85d[23] = data_0n[23];
  assign read_85d[24] = data_0n[24];
  assign read_85d[25] = data_0n[25];
  assign read_85d[26] = data_0n[26];
  assign read_85d[27] = data_0n[27];
  assign read_85d[28] = data_0n[28];
  assign read_85d[29] = data_0n[29];
  assign read_85d[30] = data_0n[30];
  assign read_85d[31] = data_0n[31];
  assign read_85d[32] = data_0n[32];
  assign read_84d[0] = data_0n[0];
  assign read_84d[1] = data_0n[1];
  assign read_84d[2] = data_0n[2];
  assign read_84d[3] = data_0n[3];
  assign read_84d[4] = data_0n[4];
  assign read_84d[5] = data_0n[5];
  assign read_84d[6] = data_0n[6];
  assign read_84d[7] = data_0n[7];
  assign read_84d[8] = data_0n[8];
  assign read_84d[9] = data_0n[9];
  assign read_84d[10] = data_0n[10];
  assign read_84d[11] = data_0n[11];
  assign read_84d[12] = data_0n[12];
  assign read_84d[13] = data_0n[13];
  assign read_84d[14] = data_0n[14];
  assign read_84d[15] = data_0n[15];
  assign read_84d[16] = data_0n[16];
  assign read_84d[17] = data_0n[17];
  assign read_84d[18] = data_0n[18];
  assign read_84d[19] = data_0n[19];
  assign read_84d[20] = data_0n[20];
  assign read_84d[21] = data_0n[21];
  assign read_84d[22] = data_0n[22];
  assign read_84d[23] = data_0n[23];
  assign read_84d[24] = data_0n[24];
  assign read_84d[25] = data_0n[25];
  assign read_84d[26] = data_0n[26];
  assign read_84d[27] = data_0n[27];
  assign read_84d[28] = data_0n[28];
  assign read_84d[29] = data_0n[29];
  assign read_84d[30] = data_0n[30];
  assign read_84d[31] = data_0n[31];
  assign read_84d[32] = data_0n[32];
  assign read_83d = data_0n[0];
  assign read_82d = data_0n[1];
  assign read_81d = data_0n[0];
  assign read_80d = data_0n[1];
  assign read_79d = data_0n[32];
  assign read_78d[0] = data_0n[1];
  assign read_78d[1] = data_0n[2];
  assign read_78d[2] = data_0n[3];
  assign read_78d[3] = data_0n[4];
  assign read_78d[4] = data_0n[5];
  assign read_78d[5] = data_0n[6];
  assign read_78d[6] = data_0n[7];
  assign read_78d[7] = data_0n[8];
  assign read_78d[8] = data_0n[9];
  assign read_78d[9] = data_0n[10];
  assign read_78d[10] = data_0n[11];
  assign read_78d[11] = data_0n[12];
  assign read_78d[12] = data_0n[13];
  assign read_78d[13] = data_0n[14];
  assign read_78d[14] = data_0n[15];
  assign read_78d[15] = data_0n[16];
  assign read_78d[16] = data_0n[17];
  assign read_78d[17] = data_0n[18];
  assign read_78d[18] = data_0n[19];
  assign read_78d[19] = data_0n[20];
  assign read_78d[20] = data_0n[21];
  assign read_78d[21] = data_0n[22];
  assign read_78d[22] = data_0n[23];
  assign read_78d[23] = data_0n[24];
  assign read_78d[24] = data_0n[25];
  assign read_78d[25] = data_0n[26];
  assign read_78d[26] = data_0n[27];
  assign read_78d[27] = data_0n[28];
  assign read_78d[28] = data_0n[29];
  assign read_78d[29] = data_0n[30];
  assign read_78d[30] = data_0n[31];
  assign read_78d[31] = data_0n[32];
  assign read_77d[0] = data_0n[0];
  assign read_77d[1] = data_0n[1];
  assign read_77d[2] = data_0n[2];
  assign read_77d[3] = data_0n[3];
  assign read_77d[4] = data_0n[4];
  assign read_77d[5] = data_0n[5];
  assign read_77d[6] = data_0n[6];
  assign read_77d[7] = data_0n[7];
  assign read_77d[8] = data_0n[8];
  assign read_77d[9] = data_0n[9];
  assign read_77d[10] = data_0n[10];
  assign read_77d[11] = data_0n[11];
  assign read_77d[12] = data_0n[12];
  assign read_77d[13] = data_0n[13];
  assign read_77d[14] = data_0n[14];
  assign read_77d[15] = data_0n[15];
  assign read_77d[16] = data_0n[16];
  assign read_77d[17] = data_0n[17];
  assign read_77d[18] = data_0n[18];
  assign read_77d[19] = data_0n[19];
  assign read_77d[20] = data_0n[20];
  assign read_77d[21] = data_0n[21];
  assign read_77d[22] = data_0n[22];
  assign read_77d[23] = data_0n[23];
  assign read_77d[24] = data_0n[24];
  assign read_77d[25] = data_0n[25];
  assign read_77d[26] = data_0n[26];
  assign read_77d[27] = data_0n[27];
  assign read_77d[28] = data_0n[28];
  assign read_77d[29] = data_0n[29];
  assign read_77d[30] = data_0n[30];
  assign read_77d[31] = data_0n[31];
  assign read_77d[32] = data_0n[32];
  assign read_76d[0] = data_0n[0];
  assign read_76d[1] = data_0n[1];
  assign read_76d[2] = data_0n[2];
  assign read_76d[3] = data_0n[3];
  assign read_76d[4] = data_0n[4];
  assign read_76d[5] = data_0n[5];
  assign read_76d[6] = data_0n[6];
  assign read_76d[7] = data_0n[7];
  assign read_76d[8] = data_0n[8];
  assign read_76d[9] = data_0n[9];
  assign read_76d[10] = data_0n[10];
  assign read_76d[11] = data_0n[11];
  assign read_76d[12] = data_0n[12];
  assign read_76d[13] = data_0n[13];
  assign read_76d[14] = data_0n[14];
  assign read_76d[15] = data_0n[15];
  assign read_76d[16] = data_0n[16];
  assign read_76d[17] = data_0n[17];
  assign read_76d[18] = data_0n[18];
  assign read_76d[19] = data_0n[19];
  assign read_76d[20] = data_0n[20];
  assign read_76d[21] = data_0n[21];
  assign read_76d[22] = data_0n[22];
  assign read_76d[23] = data_0n[23];
  assign read_76d[24] = data_0n[24];
  assign read_76d[25] = data_0n[25];
  assign read_76d[26] = data_0n[26];
  assign read_76d[27] = data_0n[27];
  assign read_76d[28] = data_0n[28];
  assign read_76d[29] = data_0n[29];
  assign read_76d[30] = data_0n[30];
  assign read_76d[31] = data_0n[31];
  assign read_76d[32] = data_0n[32];
  assign read_75d[0] = data_0n[0];
  assign read_75d[1] = data_0n[1];
  assign read_75d[2] = data_0n[2];
  assign read_75d[3] = data_0n[3];
  assign read_75d[4] = data_0n[4];
  assign read_75d[5] = data_0n[5];
  assign read_75d[6] = data_0n[6];
  assign read_75d[7] = data_0n[7];
  assign read_75d[8] = data_0n[8];
  assign read_75d[9] = data_0n[9];
  assign read_75d[10] = data_0n[10];
  assign read_75d[11] = data_0n[11];
  assign read_75d[12] = data_0n[12];
  assign read_75d[13] = data_0n[13];
  assign read_75d[14] = data_0n[14];
  assign read_75d[15] = data_0n[15];
  assign read_75d[16] = data_0n[16];
  assign read_75d[17] = data_0n[17];
  assign read_75d[18] = data_0n[18];
  assign read_75d[19] = data_0n[19];
  assign read_75d[20] = data_0n[20];
  assign read_75d[21] = data_0n[21];
  assign read_75d[22] = data_0n[22];
  assign read_75d[23] = data_0n[23];
  assign read_75d[24] = data_0n[24];
  assign read_75d[25] = data_0n[25];
  assign read_75d[26] = data_0n[26];
  assign read_75d[27] = data_0n[27];
  assign read_75d[28] = data_0n[28];
  assign read_75d[29] = data_0n[29];
  assign read_75d[30] = data_0n[30];
  assign read_75d[31] = data_0n[31];
  assign read_75d[32] = data_0n[32];
  assign read_74d[0] = data_0n[0];
  assign read_74d[1] = data_0n[1];
  assign read_74d[2] = data_0n[2];
  assign read_74d[3] = data_0n[3];
  assign read_74d[4] = data_0n[4];
  assign read_74d[5] = data_0n[5];
  assign read_74d[6] = data_0n[6];
  assign read_74d[7] = data_0n[7];
  assign read_74d[8] = data_0n[8];
  assign read_74d[9] = data_0n[9];
  assign read_74d[10] = data_0n[10];
  assign read_74d[11] = data_0n[11];
  assign read_74d[12] = data_0n[12];
  assign read_74d[13] = data_0n[13];
  assign read_74d[14] = data_0n[14];
  assign read_74d[15] = data_0n[15];
  assign read_74d[16] = data_0n[16];
  assign read_74d[17] = data_0n[17];
  assign read_74d[18] = data_0n[18];
  assign read_74d[19] = data_0n[19];
  assign read_74d[20] = data_0n[20];
  assign read_74d[21] = data_0n[21];
  assign read_74d[22] = data_0n[22];
  assign read_74d[23] = data_0n[23];
  assign read_74d[24] = data_0n[24];
  assign read_74d[25] = data_0n[25];
  assign read_74d[26] = data_0n[26];
  assign read_74d[27] = data_0n[27];
  assign read_74d[28] = data_0n[28];
  assign read_74d[29] = data_0n[29];
  assign read_74d[30] = data_0n[30];
  assign read_74d[31] = data_0n[31];
  assign read_74d[32] = data_0n[32];
  assign read_73d = data_0n[0];
  assign read_72d = data_0n[1];
  assign read_71d = data_0n[0];
  assign read_70d = data_0n[1];
  assign read_69d = data_0n[32];
  assign read_68d[0] = data_0n[1];
  assign read_68d[1] = data_0n[2];
  assign read_68d[2] = data_0n[3];
  assign read_68d[3] = data_0n[4];
  assign read_68d[4] = data_0n[5];
  assign read_68d[5] = data_0n[6];
  assign read_68d[6] = data_0n[7];
  assign read_68d[7] = data_0n[8];
  assign read_68d[8] = data_0n[9];
  assign read_68d[9] = data_0n[10];
  assign read_68d[10] = data_0n[11];
  assign read_68d[11] = data_0n[12];
  assign read_68d[12] = data_0n[13];
  assign read_68d[13] = data_0n[14];
  assign read_68d[14] = data_0n[15];
  assign read_68d[15] = data_0n[16];
  assign read_68d[16] = data_0n[17];
  assign read_68d[17] = data_0n[18];
  assign read_68d[18] = data_0n[19];
  assign read_68d[19] = data_0n[20];
  assign read_68d[20] = data_0n[21];
  assign read_68d[21] = data_0n[22];
  assign read_68d[22] = data_0n[23];
  assign read_68d[23] = data_0n[24];
  assign read_68d[24] = data_0n[25];
  assign read_68d[25] = data_0n[26];
  assign read_68d[26] = data_0n[27];
  assign read_68d[27] = data_0n[28];
  assign read_68d[28] = data_0n[29];
  assign read_68d[29] = data_0n[30];
  assign read_68d[30] = data_0n[31];
  assign read_68d[31] = data_0n[32];
  assign read_67d[0] = data_0n[0];
  assign read_67d[1] = data_0n[1];
  assign read_67d[2] = data_0n[2];
  assign read_67d[3] = data_0n[3];
  assign read_67d[4] = data_0n[4];
  assign read_67d[5] = data_0n[5];
  assign read_67d[6] = data_0n[6];
  assign read_67d[7] = data_0n[7];
  assign read_67d[8] = data_0n[8];
  assign read_67d[9] = data_0n[9];
  assign read_67d[10] = data_0n[10];
  assign read_67d[11] = data_0n[11];
  assign read_67d[12] = data_0n[12];
  assign read_67d[13] = data_0n[13];
  assign read_67d[14] = data_0n[14];
  assign read_67d[15] = data_0n[15];
  assign read_67d[16] = data_0n[16];
  assign read_67d[17] = data_0n[17];
  assign read_67d[18] = data_0n[18];
  assign read_67d[19] = data_0n[19];
  assign read_67d[20] = data_0n[20];
  assign read_67d[21] = data_0n[21];
  assign read_67d[22] = data_0n[22];
  assign read_67d[23] = data_0n[23];
  assign read_67d[24] = data_0n[24];
  assign read_67d[25] = data_0n[25];
  assign read_67d[26] = data_0n[26];
  assign read_67d[27] = data_0n[27];
  assign read_67d[28] = data_0n[28];
  assign read_67d[29] = data_0n[29];
  assign read_67d[30] = data_0n[30];
  assign read_67d[31] = data_0n[31];
  assign read_67d[32] = data_0n[32];
  assign read_66d[0] = data_0n[0];
  assign read_66d[1] = data_0n[1];
  assign read_66d[2] = data_0n[2];
  assign read_66d[3] = data_0n[3];
  assign read_66d[4] = data_0n[4];
  assign read_66d[5] = data_0n[5];
  assign read_66d[6] = data_0n[6];
  assign read_66d[7] = data_0n[7];
  assign read_66d[8] = data_0n[8];
  assign read_66d[9] = data_0n[9];
  assign read_66d[10] = data_0n[10];
  assign read_66d[11] = data_0n[11];
  assign read_66d[12] = data_0n[12];
  assign read_66d[13] = data_0n[13];
  assign read_66d[14] = data_0n[14];
  assign read_66d[15] = data_0n[15];
  assign read_66d[16] = data_0n[16];
  assign read_66d[17] = data_0n[17];
  assign read_66d[18] = data_0n[18];
  assign read_66d[19] = data_0n[19];
  assign read_66d[20] = data_0n[20];
  assign read_66d[21] = data_0n[21];
  assign read_66d[22] = data_0n[22];
  assign read_66d[23] = data_0n[23];
  assign read_66d[24] = data_0n[24];
  assign read_66d[25] = data_0n[25];
  assign read_66d[26] = data_0n[26];
  assign read_66d[27] = data_0n[27];
  assign read_66d[28] = data_0n[28];
  assign read_66d[29] = data_0n[29];
  assign read_66d[30] = data_0n[30];
  assign read_66d[31] = data_0n[31];
  assign read_66d[32] = data_0n[32];
  assign read_65d[0] = data_0n[0];
  assign read_65d[1] = data_0n[1];
  assign read_65d[2] = data_0n[2];
  assign read_65d[3] = data_0n[3];
  assign read_65d[4] = data_0n[4];
  assign read_65d[5] = data_0n[5];
  assign read_65d[6] = data_0n[6];
  assign read_65d[7] = data_0n[7];
  assign read_65d[8] = data_0n[8];
  assign read_65d[9] = data_0n[9];
  assign read_65d[10] = data_0n[10];
  assign read_65d[11] = data_0n[11];
  assign read_65d[12] = data_0n[12];
  assign read_65d[13] = data_0n[13];
  assign read_65d[14] = data_0n[14];
  assign read_65d[15] = data_0n[15];
  assign read_65d[16] = data_0n[16];
  assign read_65d[17] = data_0n[17];
  assign read_65d[18] = data_0n[18];
  assign read_65d[19] = data_0n[19];
  assign read_65d[20] = data_0n[20];
  assign read_65d[21] = data_0n[21];
  assign read_65d[22] = data_0n[22];
  assign read_65d[23] = data_0n[23];
  assign read_65d[24] = data_0n[24];
  assign read_65d[25] = data_0n[25];
  assign read_65d[26] = data_0n[26];
  assign read_65d[27] = data_0n[27];
  assign read_65d[28] = data_0n[28];
  assign read_65d[29] = data_0n[29];
  assign read_65d[30] = data_0n[30];
  assign read_65d[31] = data_0n[31];
  assign read_65d[32] = data_0n[32];
  assign read_64d[0] = data_0n[0];
  assign read_64d[1] = data_0n[1];
  assign read_64d[2] = data_0n[2];
  assign read_64d[3] = data_0n[3];
  assign read_64d[4] = data_0n[4];
  assign read_64d[5] = data_0n[5];
  assign read_64d[6] = data_0n[6];
  assign read_64d[7] = data_0n[7];
  assign read_64d[8] = data_0n[8];
  assign read_64d[9] = data_0n[9];
  assign read_64d[10] = data_0n[10];
  assign read_64d[11] = data_0n[11];
  assign read_64d[12] = data_0n[12];
  assign read_64d[13] = data_0n[13];
  assign read_64d[14] = data_0n[14];
  assign read_64d[15] = data_0n[15];
  assign read_64d[16] = data_0n[16];
  assign read_64d[17] = data_0n[17];
  assign read_64d[18] = data_0n[18];
  assign read_64d[19] = data_0n[19];
  assign read_64d[20] = data_0n[20];
  assign read_64d[21] = data_0n[21];
  assign read_64d[22] = data_0n[22];
  assign read_64d[23] = data_0n[23];
  assign read_64d[24] = data_0n[24];
  assign read_64d[25] = data_0n[25];
  assign read_64d[26] = data_0n[26];
  assign read_64d[27] = data_0n[27];
  assign read_64d[28] = data_0n[28];
  assign read_64d[29] = data_0n[29];
  assign read_64d[30] = data_0n[30];
  assign read_64d[31] = data_0n[31];
  assign read_64d[32] = data_0n[32];
  assign read_63d = data_0n[0];
  assign read_62d = data_0n[1];
  assign read_61d = data_0n[0];
  assign read_60d = data_0n[1];
  assign read_59d = data_0n[32];
  assign read_58d[0] = data_0n[1];
  assign read_58d[1] = data_0n[2];
  assign read_58d[2] = data_0n[3];
  assign read_58d[3] = data_0n[4];
  assign read_58d[4] = data_0n[5];
  assign read_58d[5] = data_0n[6];
  assign read_58d[6] = data_0n[7];
  assign read_58d[7] = data_0n[8];
  assign read_58d[8] = data_0n[9];
  assign read_58d[9] = data_0n[10];
  assign read_58d[10] = data_0n[11];
  assign read_58d[11] = data_0n[12];
  assign read_58d[12] = data_0n[13];
  assign read_58d[13] = data_0n[14];
  assign read_58d[14] = data_0n[15];
  assign read_58d[15] = data_0n[16];
  assign read_58d[16] = data_0n[17];
  assign read_58d[17] = data_0n[18];
  assign read_58d[18] = data_0n[19];
  assign read_58d[19] = data_0n[20];
  assign read_58d[20] = data_0n[21];
  assign read_58d[21] = data_0n[22];
  assign read_58d[22] = data_0n[23];
  assign read_58d[23] = data_0n[24];
  assign read_58d[24] = data_0n[25];
  assign read_58d[25] = data_0n[26];
  assign read_58d[26] = data_0n[27];
  assign read_58d[27] = data_0n[28];
  assign read_58d[28] = data_0n[29];
  assign read_58d[29] = data_0n[30];
  assign read_58d[30] = data_0n[31];
  assign read_58d[31] = data_0n[32];
  assign read_57d[0] = data_0n[0];
  assign read_57d[1] = data_0n[1];
  assign read_57d[2] = data_0n[2];
  assign read_57d[3] = data_0n[3];
  assign read_57d[4] = data_0n[4];
  assign read_57d[5] = data_0n[5];
  assign read_57d[6] = data_0n[6];
  assign read_57d[7] = data_0n[7];
  assign read_57d[8] = data_0n[8];
  assign read_57d[9] = data_0n[9];
  assign read_57d[10] = data_0n[10];
  assign read_57d[11] = data_0n[11];
  assign read_57d[12] = data_0n[12];
  assign read_57d[13] = data_0n[13];
  assign read_57d[14] = data_0n[14];
  assign read_57d[15] = data_0n[15];
  assign read_57d[16] = data_0n[16];
  assign read_57d[17] = data_0n[17];
  assign read_57d[18] = data_0n[18];
  assign read_57d[19] = data_0n[19];
  assign read_57d[20] = data_0n[20];
  assign read_57d[21] = data_0n[21];
  assign read_57d[22] = data_0n[22];
  assign read_57d[23] = data_0n[23];
  assign read_57d[24] = data_0n[24];
  assign read_57d[25] = data_0n[25];
  assign read_57d[26] = data_0n[26];
  assign read_57d[27] = data_0n[27];
  assign read_57d[28] = data_0n[28];
  assign read_57d[29] = data_0n[29];
  assign read_57d[30] = data_0n[30];
  assign read_57d[31] = data_0n[31];
  assign read_57d[32] = data_0n[32];
  assign read_56d[0] = data_0n[0];
  assign read_56d[1] = data_0n[1];
  assign read_56d[2] = data_0n[2];
  assign read_56d[3] = data_0n[3];
  assign read_56d[4] = data_0n[4];
  assign read_56d[5] = data_0n[5];
  assign read_56d[6] = data_0n[6];
  assign read_56d[7] = data_0n[7];
  assign read_56d[8] = data_0n[8];
  assign read_56d[9] = data_0n[9];
  assign read_56d[10] = data_0n[10];
  assign read_56d[11] = data_0n[11];
  assign read_56d[12] = data_0n[12];
  assign read_56d[13] = data_0n[13];
  assign read_56d[14] = data_0n[14];
  assign read_56d[15] = data_0n[15];
  assign read_56d[16] = data_0n[16];
  assign read_56d[17] = data_0n[17];
  assign read_56d[18] = data_0n[18];
  assign read_56d[19] = data_0n[19];
  assign read_56d[20] = data_0n[20];
  assign read_56d[21] = data_0n[21];
  assign read_56d[22] = data_0n[22];
  assign read_56d[23] = data_0n[23];
  assign read_56d[24] = data_0n[24];
  assign read_56d[25] = data_0n[25];
  assign read_56d[26] = data_0n[26];
  assign read_56d[27] = data_0n[27];
  assign read_56d[28] = data_0n[28];
  assign read_56d[29] = data_0n[29];
  assign read_56d[30] = data_0n[30];
  assign read_56d[31] = data_0n[31];
  assign read_56d[32] = data_0n[32];
  assign read_55d[0] = data_0n[0];
  assign read_55d[1] = data_0n[1];
  assign read_55d[2] = data_0n[2];
  assign read_55d[3] = data_0n[3];
  assign read_55d[4] = data_0n[4];
  assign read_55d[5] = data_0n[5];
  assign read_55d[6] = data_0n[6];
  assign read_55d[7] = data_0n[7];
  assign read_55d[8] = data_0n[8];
  assign read_55d[9] = data_0n[9];
  assign read_55d[10] = data_0n[10];
  assign read_55d[11] = data_0n[11];
  assign read_55d[12] = data_0n[12];
  assign read_55d[13] = data_0n[13];
  assign read_55d[14] = data_0n[14];
  assign read_55d[15] = data_0n[15];
  assign read_55d[16] = data_0n[16];
  assign read_55d[17] = data_0n[17];
  assign read_55d[18] = data_0n[18];
  assign read_55d[19] = data_0n[19];
  assign read_55d[20] = data_0n[20];
  assign read_55d[21] = data_0n[21];
  assign read_55d[22] = data_0n[22];
  assign read_55d[23] = data_0n[23];
  assign read_55d[24] = data_0n[24];
  assign read_55d[25] = data_0n[25];
  assign read_55d[26] = data_0n[26];
  assign read_55d[27] = data_0n[27];
  assign read_55d[28] = data_0n[28];
  assign read_55d[29] = data_0n[29];
  assign read_55d[30] = data_0n[30];
  assign read_55d[31] = data_0n[31];
  assign read_55d[32] = data_0n[32];
  assign read_54d[0] = data_0n[0];
  assign read_54d[1] = data_0n[1];
  assign read_54d[2] = data_0n[2];
  assign read_54d[3] = data_0n[3];
  assign read_54d[4] = data_0n[4];
  assign read_54d[5] = data_0n[5];
  assign read_54d[6] = data_0n[6];
  assign read_54d[7] = data_0n[7];
  assign read_54d[8] = data_0n[8];
  assign read_54d[9] = data_0n[9];
  assign read_54d[10] = data_0n[10];
  assign read_54d[11] = data_0n[11];
  assign read_54d[12] = data_0n[12];
  assign read_54d[13] = data_0n[13];
  assign read_54d[14] = data_0n[14];
  assign read_54d[15] = data_0n[15];
  assign read_54d[16] = data_0n[16];
  assign read_54d[17] = data_0n[17];
  assign read_54d[18] = data_0n[18];
  assign read_54d[19] = data_0n[19];
  assign read_54d[20] = data_0n[20];
  assign read_54d[21] = data_0n[21];
  assign read_54d[22] = data_0n[22];
  assign read_54d[23] = data_0n[23];
  assign read_54d[24] = data_0n[24];
  assign read_54d[25] = data_0n[25];
  assign read_54d[26] = data_0n[26];
  assign read_54d[27] = data_0n[27];
  assign read_54d[28] = data_0n[28];
  assign read_54d[29] = data_0n[29];
  assign read_54d[30] = data_0n[30];
  assign read_54d[31] = data_0n[31];
  assign read_54d[32] = data_0n[32];
  assign read_53d = data_0n[0];
  assign read_52d = data_0n[1];
  assign read_51d = data_0n[0];
  assign read_50d = data_0n[1];
  assign read_49d = data_0n[32];
  assign read_48d[0] = data_0n[1];
  assign read_48d[1] = data_0n[2];
  assign read_48d[2] = data_0n[3];
  assign read_48d[3] = data_0n[4];
  assign read_48d[4] = data_0n[5];
  assign read_48d[5] = data_0n[6];
  assign read_48d[6] = data_0n[7];
  assign read_48d[7] = data_0n[8];
  assign read_48d[8] = data_0n[9];
  assign read_48d[9] = data_0n[10];
  assign read_48d[10] = data_0n[11];
  assign read_48d[11] = data_0n[12];
  assign read_48d[12] = data_0n[13];
  assign read_48d[13] = data_0n[14];
  assign read_48d[14] = data_0n[15];
  assign read_48d[15] = data_0n[16];
  assign read_48d[16] = data_0n[17];
  assign read_48d[17] = data_0n[18];
  assign read_48d[18] = data_0n[19];
  assign read_48d[19] = data_0n[20];
  assign read_48d[20] = data_0n[21];
  assign read_48d[21] = data_0n[22];
  assign read_48d[22] = data_0n[23];
  assign read_48d[23] = data_0n[24];
  assign read_48d[24] = data_0n[25];
  assign read_48d[25] = data_0n[26];
  assign read_48d[26] = data_0n[27];
  assign read_48d[27] = data_0n[28];
  assign read_48d[28] = data_0n[29];
  assign read_48d[29] = data_0n[30];
  assign read_48d[30] = data_0n[31];
  assign read_48d[31] = data_0n[32];
  assign read_47d[0] = data_0n[0];
  assign read_47d[1] = data_0n[1];
  assign read_47d[2] = data_0n[2];
  assign read_47d[3] = data_0n[3];
  assign read_47d[4] = data_0n[4];
  assign read_47d[5] = data_0n[5];
  assign read_47d[6] = data_0n[6];
  assign read_47d[7] = data_0n[7];
  assign read_47d[8] = data_0n[8];
  assign read_47d[9] = data_0n[9];
  assign read_47d[10] = data_0n[10];
  assign read_47d[11] = data_0n[11];
  assign read_47d[12] = data_0n[12];
  assign read_47d[13] = data_0n[13];
  assign read_47d[14] = data_0n[14];
  assign read_47d[15] = data_0n[15];
  assign read_47d[16] = data_0n[16];
  assign read_47d[17] = data_0n[17];
  assign read_47d[18] = data_0n[18];
  assign read_47d[19] = data_0n[19];
  assign read_47d[20] = data_0n[20];
  assign read_47d[21] = data_0n[21];
  assign read_47d[22] = data_0n[22];
  assign read_47d[23] = data_0n[23];
  assign read_47d[24] = data_0n[24];
  assign read_47d[25] = data_0n[25];
  assign read_47d[26] = data_0n[26];
  assign read_47d[27] = data_0n[27];
  assign read_47d[28] = data_0n[28];
  assign read_47d[29] = data_0n[29];
  assign read_47d[30] = data_0n[30];
  assign read_47d[31] = data_0n[31];
  assign read_47d[32] = data_0n[32];
  assign read_46d[0] = data_0n[0];
  assign read_46d[1] = data_0n[1];
  assign read_46d[2] = data_0n[2];
  assign read_46d[3] = data_0n[3];
  assign read_46d[4] = data_0n[4];
  assign read_46d[5] = data_0n[5];
  assign read_46d[6] = data_0n[6];
  assign read_46d[7] = data_0n[7];
  assign read_46d[8] = data_0n[8];
  assign read_46d[9] = data_0n[9];
  assign read_46d[10] = data_0n[10];
  assign read_46d[11] = data_0n[11];
  assign read_46d[12] = data_0n[12];
  assign read_46d[13] = data_0n[13];
  assign read_46d[14] = data_0n[14];
  assign read_46d[15] = data_0n[15];
  assign read_46d[16] = data_0n[16];
  assign read_46d[17] = data_0n[17];
  assign read_46d[18] = data_0n[18];
  assign read_46d[19] = data_0n[19];
  assign read_46d[20] = data_0n[20];
  assign read_46d[21] = data_0n[21];
  assign read_46d[22] = data_0n[22];
  assign read_46d[23] = data_0n[23];
  assign read_46d[24] = data_0n[24];
  assign read_46d[25] = data_0n[25];
  assign read_46d[26] = data_0n[26];
  assign read_46d[27] = data_0n[27];
  assign read_46d[28] = data_0n[28];
  assign read_46d[29] = data_0n[29];
  assign read_46d[30] = data_0n[30];
  assign read_46d[31] = data_0n[31];
  assign read_46d[32] = data_0n[32];
  assign read_45d[0] = data_0n[0];
  assign read_45d[1] = data_0n[1];
  assign read_45d[2] = data_0n[2];
  assign read_45d[3] = data_0n[3];
  assign read_45d[4] = data_0n[4];
  assign read_45d[5] = data_0n[5];
  assign read_45d[6] = data_0n[6];
  assign read_45d[7] = data_0n[7];
  assign read_45d[8] = data_0n[8];
  assign read_45d[9] = data_0n[9];
  assign read_45d[10] = data_0n[10];
  assign read_45d[11] = data_0n[11];
  assign read_45d[12] = data_0n[12];
  assign read_45d[13] = data_0n[13];
  assign read_45d[14] = data_0n[14];
  assign read_45d[15] = data_0n[15];
  assign read_45d[16] = data_0n[16];
  assign read_45d[17] = data_0n[17];
  assign read_45d[18] = data_0n[18];
  assign read_45d[19] = data_0n[19];
  assign read_45d[20] = data_0n[20];
  assign read_45d[21] = data_0n[21];
  assign read_45d[22] = data_0n[22];
  assign read_45d[23] = data_0n[23];
  assign read_45d[24] = data_0n[24];
  assign read_45d[25] = data_0n[25];
  assign read_45d[26] = data_0n[26];
  assign read_45d[27] = data_0n[27];
  assign read_45d[28] = data_0n[28];
  assign read_45d[29] = data_0n[29];
  assign read_45d[30] = data_0n[30];
  assign read_45d[31] = data_0n[31];
  assign read_45d[32] = data_0n[32];
  assign read_44d[0] = data_0n[0];
  assign read_44d[1] = data_0n[1];
  assign read_44d[2] = data_0n[2];
  assign read_44d[3] = data_0n[3];
  assign read_44d[4] = data_0n[4];
  assign read_44d[5] = data_0n[5];
  assign read_44d[6] = data_0n[6];
  assign read_44d[7] = data_0n[7];
  assign read_44d[8] = data_0n[8];
  assign read_44d[9] = data_0n[9];
  assign read_44d[10] = data_0n[10];
  assign read_44d[11] = data_0n[11];
  assign read_44d[12] = data_0n[12];
  assign read_44d[13] = data_0n[13];
  assign read_44d[14] = data_0n[14];
  assign read_44d[15] = data_0n[15];
  assign read_44d[16] = data_0n[16];
  assign read_44d[17] = data_0n[17];
  assign read_44d[18] = data_0n[18];
  assign read_44d[19] = data_0n[19];
  assign read_44d[20] = data_0n[20];
  assign read_44d[21] = data_0n[21];
  assign read_44d[22] = data_0n[22];
  assign read_44d[23] = data_0n[23];
  assign read_44d[24] = data_0n[24];
  assign read_44d[25] = data_0n[25];
  assign read_44d[26] = data_0n[26];
  assign read_44d[27] = data_0n[27];
  assign read_44d[28] = data_0n[28];
  assign read_44d[29] = data_0n[29];
  assign read_44d[30] = data_0n[30];
  assign read_44d[31] = data_0n[31];
  assign read_44d[32] = data_0n[32];
  assign read_43d = data_0n[0];
  assign read_42d = data_0n[1];
  assign read_41d = data_0n[0];
  assign read_40d = data_0n[1];
  assign read_39d = data_0n[32];
  assign read_38d[0] = data_0n[1];
  assign read_38d[1] = data_0n[2];
  assign read_38d[2] = data_0n[3];
  assign read_38d[3] = data_0n[4];
  assign read_38d[4] = data_0n[5];
  assign read_38d[5] = data_0n[6];
  assign read_38d[6] = data_0n[7];
  assign read_38d[7] = data_0n[8];
  assign read_38d[8] = data_0n[9];
  assign read_38d[9] = data_0n[10];
  assign read_38d[10] = data_0n[11];
  assign read_38d[11] = data_0n[12];
  assign read_38d[12] = data_0n[13];
  assign read_38d[13] = data_0n[14];
  assign read_38d[14] = data_0n[15];
  assign read_38d[15] = data_0n[16];
  assign read_38d[16] = data_0n[17];
  assign read_38d[17] = data_0n[18];
  assign read_38d[18] = data_0n[19];
  assign read_38d[19] = data_0n[20];
  assign read_38d[20] = data_0n[21];
  assign read_38d[21] = data_0n[22];
  assign read_38d[22] = data_0n[23];
  assign read_38d[23] = data_0n[24];
  assign read_38d[24] = data_0n[25];
  assign read_38d[25] = data_0n[26];
  assign read_38d[26] = data_0n[27];
  assign read_38d[27] = data_0n[28];
  assign read_38d[28] = data_0n[29];
  assign read_38d[29] = data_0n[30];
  assign read_38d[30] = data_0n[31];
  assign read_38d[31] = data_0n[32];
  assign read_37d[0] = data_0n[0];
  assign read_37d[1] = data_0n[1];
  assign read_37d[2] = data_0n[2];
  assign read_37d[3] = data_0n[3];
  assign read_37d[4] = data_0n[4];
  assign read_37d[5] = data_0n[5];
  assign read_37d[6] = data_0n[6];
  assign read_37d[7] = data_0n[7];
  assign read_37d[8] = data_0n[8];
  assign read_37d[9] = data_0n[9];
  assign read_37d[10] = data_0n[10];
  assign read_37d[11] = data_0n[11];
  assign read_37d[12] = data_0n[12];
  assign read_37d[13] = data_0n[13];
  assign read_37d[14] = data_0n[14];
  assign read_37d[15] = data_0n[15];
  assign read_37d[16] = data_0n[16];
  assign read_37d[17] = data_0n[17];
  assign read_37d[18] = data_0n[18];
  assign read_37d[19] = data_0n[19];
  assign read_37d[20] = data_0n[20];
  assign read_37d[21] = data_0n[21];
  assign read_37d[22] = data_0n[22];
  assign read_37d[23] = data_0n[23];
  assign read_37d[24] = data_0n[24];
  assign read_37d[25] = data_0n[25];
  assign read_37d[26] = data_0n[26];
  assign read_37d[27] = data_0n[27];
  assign read_37d[28] = data_0n[28];
  assign read_37d[29] = data_0n[29];
  assign read_37d[30] = data_0n[30];
  assign read_37d[31] = data_0n[31];
  assign read_37d[32] = data_0n[32];
  assign read_36d[0] = data_0n[0];
  assign read_36d[1] = data_0n[1];
  assign read_36d[2] = data_0n[2];
  assign read_36d[3] = data_0n[3];
  assign read_36d[4] = data_0n[4];
  assign read_36d[5] = data_0n[5];
  assign read_36d[6] = data_0n[6];
  assign read_36d[7] = data_0n[7];
  assign read_36d[8] = data_0n[8];
  assign read_36d[9] = data_0n[9];
  assign read_36d[10] = data_0n[10];
  assign read_36d[11] = data_0n[11];
  assign read_36d[12] = data_0n[12];
  assign read_36d[13] = data_0n[13];
  assign read_36d[14] = data_0n[14];
  assign read_36d[15] = data_0n[15];
  assign read_36d[16] = data_0n[16];
  assign read_36d[17] = data_0n[17];
  assign read_36d[18] = data_0n[18];
  assign read_36d[19] = data_0n[19];
  assign read_36d[20] = data_0n[20];
  assign read_36d[21] = data_0n[21];
  assign read_36d[22] = data_0n[22];
  assign read_36d[23] = data_0n[23];
  assign read_36d[24] = data_0n[24];
  assign read_36d[25] = data_0n[25];
  assign read_36d[26] = data_0n[26];
  assign read_36d[27] = data_0n[27];
  assign read_36d[28] = data_0n[28];
  assign read_36d[29] = data_0n[29];
  assign read_36d[30] = data_0n[30];
  assign read_36d[31] = data_0n[31];
  assign read_36d[32] = data_0n[32];
  assign read_35d[0] = data_0n[0];
  assign read_35d[1] = data_0n[1];
  assign read_35d[2] = data_0n[2];
  assign read_35d[3] = data_0n[3];
  assign read_35d[4] = data_0n[4];
  assign read_35d[5] = data_0n[5];
  assign read_35d[6] = data_0n[6];
  assign read_35d[7] = data_0n[7];
  assign read_35d[8] = data_0n[8];
  assign read_35d[9] = data_0n[9];
  assign read_35d[10] = data_0n[10];
  assign read_35d[11] = data_0n[11];
  assign read_35d[12] = data_0n[12];
  assign read_35d[13] = data_0n[13];
  assign read_35d[14] = data_0n[14];
  assign read_35d[15] = data_0n[15];
  assign read_35d[16] = data_0n[16];
  assign read_35d[17] = data_0n[17];
  assign read_35d[18] = data_0n[18];
  assign read_35d[19] = data_0n[19];
  assign read_35d[20] = data_0n[20];
  assign read_35d[21] = data_0n[21];
  assign read_35d[22] = data_0n[22];
  assign read_35d[23] = data_0n[23];
  assign read_35d[24] = data_0n[24];
  assign read_35d[25] = data_0n[25];
  assign read_35d[26] = data_0n[26];
  assign read_35d[27] = data_0n[27];
  assign read_35d[28] = data_0n[28];
  assign read_35d[29] = data_0n[29];
  assign read_35d[30] = data_0n[30];
  assign read_35d[31] = data_0n[31];
  assign read_35d[32] = data_0n[32];
  assign read_34d[0] = data_0n[0];
  assign read_34d[1] = data_0n[1];
  assign read_34d[2] = data_0n[2];
  assign read_34d[3] = data_0n[3];
  assign read_34d[4] = data_0n[4];
  assign read_34d[5] = data_0n[5];
  assign read_34d[6] = data_0n[6];
  assign read_34d[7] = data_0n[7];
  assign read_34d[8] = data_0n[8];
  assign read_34d[9] = data_0n[9];
  assign read_34d[10] = data_0n[10];
  assign read_34d[11] = data_0n[11];
  assign read_34d[12] = data_0n[12];
  assign read_34d[13] = data_0n[13];
  assign read_34d[14] = data_0n[14];
  assign read_34d[15] = data_0n[15];
  assign read_34d[16] = data_0n[16];
  assign read_34d[17] = data_0n[17];
  assign read_34d[18] = data_0n[18];
  assign read_34d[19] = data_0n[19];
  assign read_34d[20] = data_0n[20];
  assign read_34d[21] = data_0n[21];
  assign read_34d[22] = data_0n[22];
  assign read_34d[23] = data_0n[23];
  assign read_34d[24] = data_0n[24];
  assign read_34d[25] = data_0n[25];
  assign read_34d[26] = data_0n[26];
  assign read_34d[27] = data_0n[27];
  assign read_34d[28] = data_0n[28];
  assign read_34d[29] = data_0n[29];
  assign read_34d[30] = data_0n[30];
  assign read_34d[31] = data_0n[31];
  assign read_34d[32] = data_0n[32];
  assign read_33d = data_0n[0];
  assign read_32d = data_0n[1];
  assign read_31d = data_0n[0];
  assign read_30d = data_0n[1];
  assign read_29d = data_0n[32];
  assign read_28d[0] = data_0n[1];
  assign read_28d[1] = data_0n[2];
  assign read_28d[2] = data_0n[3];
  assign read_28d[3] = data_0n[4];
  assign read_28d[4] = data_0n[5];
  assign read_28d[5] = data_0n[6];
  assign read_28d[6] = data_0n[7];
  assign read_28d[7] = data_0n[8];
  assign read_28d[8] = data_0n[9];
  assign read_28d[9] = data_0n[10];
  assign read_28d[10] = data_0n[11];
  assign read_28d[11] = data_0n[12];
  assign read_28d[12] = data_0n[13];
  assign read_28d[13] = data_0n[14];
  assign read_28d[14] = data_0n[15];
  assign read_28d[15] = data_0n[16];
  assign read_28d[16] = data_0n[17];
  assign read_28d[17] = data_0n[18];
  assign read_28d[18] = data_0n[19];
  assign read_28d[19] = data_0n[20];
  assign read_28d[20] = data_0n[21];
  assign read_28d[21] = data_0n[22];
  assign read_28d[22] = data_0n[23];
  assign read_28d[23] = data_0n[24];
  assign read_28d[24] = data_0n[25];
  assign read_28d[25] = data_0n[26];
  assign read_28d[26] = data_0n[27];
  assign read_28d[27] = data_0n[28];
  assign read_28d[28] = data_0n[29];
  assign read_28d[29] = data_0n[30];
  assign read_28d[30] = data_0n[31];
  assign read_28d[31] = data_0n[32];
  assign read_27d[0] = data_0n[0];
  assign read_27d[1] = data_0n[1];
  assign read_27d[2] = data_0n[2];
  assign read_27d[3] = data_0n[3];
  assign read_27d[4] = data_0n[4];
  assign read_27d[5] = data_0n[5];
  assign read_27d[6] = data_0n[6];
  assign read_27d[7] = data_0n[7];
  assign read_27d[8] = data_0n[8];
  assign read_27d[9] = data_0n[9];
  assign read_27d[10] = data_0n[10];
  assign read_27d[11] = data_0n[11];
  assign read_27d[12] = data_0n[12];
  assign read_27d[13] = data_0n[13];
  assign read_27d[14] = data_0n[14];
  assign read_27d[15] = data_0n[15];
  assign read_27d[16] = data_0n[16];
  assign read_27d[17] = data_0n[17];
  assign read_27d[18] = data_0n[18];
  assign read_27d[19] = data_0n[19];
  assign read_27d[20] = data_0n[20];
  assign read_27d[21] = data_0n[21];
  assign read_27d[22] = data_0n[22];
  assign read_27d[23] = data_0n[23];
  assign read_27d[24] = data_0n[24];
  assign read_27d[25] = data_0n[25];
  assign read_27d[26] = data_0n[26];
  assign read_27d[27] = data_0n[27];
  assign read_27d[28] = data_0n[28];
  assign read_27d[29] = data_0n[29];
  assign read_27d[30] = data_0n[30];
  assign read_27d[31] = data_0n[31];
  assign read_27d[32] = data_0n[32];
  assign read_26d[0] = data_0n[0];
  assign read_26d[1] = data_0n[1];
  assign read_26d[2] = data_0n[2];
  assign read_26d[3] = data_0n[3];
  assign read_26d[4] = data_0n[4];
  assign read_26d[5] = data_0n[5];
  assign read_26d[6] = data_0n[6];
  assign read_26d[7] = data_0n[7];
  assign read_26d[8] = data_0n[8];
  assign read_26d[9] = data_0n[9];
  assign read_26d[10] = data_0n[10];
  assign read_26d[11] = data_0n[11];
  assign read_26d[12] = data_0n[12];
  assign read_26d[13] = data_0n[13];
  assign read_26d[14] = data_0n[14];
  assign read_26d[15] = data_0n[15];
  assign read_26d[16] = data_0n[16];
  assign read_26d[17] = data_0n[17];
  assign read_26d[18] = data_0n[18];
  assign read_26d[19] = data_0n[19];
  assign read_26d[20] = data_0n[20];
  assign read_26d[21] = data_0n[21];
  assign read_26d[22] = data_0n[22];
  assign read_26d[23] = data_0n[23];
  assign read_26d[24] = data_0n[24];
  assign read_26d[25] = data_0n[25];
  assign read_26d[26] = data_0n[26];
  assign read_26d[27] = data_0n[27];
  assign read_26d[28] = data_0n[28];
  assign read_26d[29] = data_0n[29];
  assign read_26d[30] = data_0n[30];
  assign read_26d[31] = data_0n[31];
  assign read_26d[32] = data_0n[32];
  assign read_25d[0] = data_0n[0];
  assign read_25d[1] = data_0n[1];
  assign read_25d[2] = data_0n[2];
  assign read_25d[3] = data_0n[3];
  assign read_25d[4] = data_0n[4];
  assign read_25d[5] = data_0n[5];
  assign read_25d[6] = data_0n[6];
  assign read_25d[7] = data_0n[7];
  assign read_25d[8] = data_0n[8];
  assign read_25d[9] = data_0n[9];
  assign read_25d[10] = data_0n[10];
  assign read_25d[11] = data_0n[11];
  assign read_25d[12] = data_0n[12];
  assign read_25d[13] = data_0n[13];
  assign read_25d[14] = data_0n[14];
  assign read_25d[15] = data_0n[15];
  assign read_25d[16] = data_0n[16];
  assign read_25d[17] = data_0n[17];
  assign read_25d[18] = data_0n[18];
  assign read_25d[19] = data_0n[19];
  assign read_25d[20] = data_0n[20];
  assign read_25d[21] = data_0n[21];
  assign read_25d[22] = data_0n[22];
  assign read_25d[23] = data_0n[23];
  assign read_25d[24] = data_0n[24];
  assign read_25d[25] = data_0n[25];
  assign read_25d[26] = data_0n[26];
  assign read_25d[27] = data_0n[27];
  assign read_25d[28] = data_0n[28];
  assign read_25d[29] = data_0n[29];
  assign read_25d[30] = data_0n[30];
  assign read_25d[31] = data_0n[31];
  assign read_25d[32] = data_0n[32];
  assign read_24d[0] = data_0n[0];
  assign read_24d[1] = data_0n[1];
  assign read_24d[2] = data_0n[2];
  assign read_24d[3] = data_0n[3];
  assign read_24d[4] = data_0n[4];
  assign read_24d[5] = data_0n[5];
  assign read_24d[6] = data_0n[6];
  assign read_24d[7] = data_0n[7];
  assign read_24d[8] = data_0n[8];
  assign read_24d[9] = data_0n[9];
  assign read_24d[10] = data_0n[10];
  assign read_24d[11] = data_0n[11];
  assign read_24d[12] = data_0n[12];
  assign read_24d[13] = data_0n[13];
  assign read_24d[14] = data_0n[14];
  assign read_24d[15] = data_0n[15];
  assign read_24d[16] = data_0n[16];
  assign read_24d[17] = data_0n[17];
  assign read_24d[18] = data_0n[18];
  assign read_24d[19] = data_0n[19];
  assign read_24d[20] = data_0n[20];
  assign read_24d[21] = data_0n[21];
  assign read_24d[22] = data_0n[22];
  assign read_24d[23] = data_0n[23];
  assign read_24d[24] = data_0n[24];
  assign read_24d[25] = data_0n[25];
  assign read_24d[26] = data_0n[26];
  assign read_24d[27] = data_0n[27];
  assign read_24d[28] = data_0n[28];
  assign read_24d[29] = data_0n[29];
  assign read_24d[30] = data_0n[30];
  assign read_24d[31] = data_0n[31];
  assign read_24d[32] = data_0n[32];
  assign read_23d = data_0n[0];
  assign read_22d = data_0n[1];
  assign read_21d = data_0n[0];
  assign read_20d = data_0n[1];
  assign read_19d = data_0n[32];
  assign read_18d[0] = data_0n[1];
  assign read_18d[1] = data_0n[2];
  assign read_18d[2] = data_0n[3];
  assign read_18d[3] = data_0n[4];
  assign read_18d[4] = data_0n[5];
  assign read_18d[5] = data_0n[6];
  assign read_18d[6] = data_0n[7];
  assign read_18d[7] = data_0n[8];
  assign read_18d[8] = data_0n[9];
  assign read_18d[9] = data_0n[10];
  assign read_18d[10] = data_0n[11];
  assign read_18d[11] = data_0n[12];
  assign read_18d[12] = data_0n[13];
  assign read_18d[13] = data_0n[14];
  assign read_18d[14] = data_0n[15];
  assign read_18d[15] = data_0n[16];
  assign read_18d[16] = data_0n[17];
  assign read_18d[17] = data_0n[18];
  assign read_18d[18] = data_0n[19];
  assign read_18d[19] = data_0n[20];
  assign read_18d[20] = data_0n[21];
  assign read_18d[21] = data_0n[22];
  assign read_18d[22] = data_0n[23];
  assign read_18d[23] = data_0n[24];
  assign read_18d[24] = data_0n[25];
  assign read_18d[25] = data_0n[26];
  assign read_18d[26] = data_0n[27];
  assign read_18d[27] = data_0n[28];
  assign read_18d[28] = data_0n[29];
  assign read_18d[29] = data_0n[30];
  assign read_18d[30] = data_0n[31];
  assign read_18d[31] = data_0n[32];
  assign read_17d[0] = data_0n[0];
  assign read_17d[1] = data_0n[1];
  assign read_17d[2] = data_0n[2];
  assign read_17d[3] = data_0n[3];
  assign read_17d[4] = data_0n[4];
  assign read_17d[5] = data_0n[5];
  assign read_17d[6] = data_0n[6];
  assign read_17d[7] = data_0n[7];
  assign read_17d[8] = data_0n[8];
  assign read_17d[9] = data_0n[9];
  assign read_17d[10] = data_0n[10];
  assign read_17d[11] = data_0n[11];
  assign read_17d[12] = data_0n[12];
  assign read_17d[13] = data_0n[13];
  assign read_17d[14] = data_0n[14];
  assign read_17d[15] = data_0n[15];
  assign read_17d[16] = data_0n[16];
  assign read_17d[17] = data_0n[17];
  assign read_17d[18] = data_0n[18];
  assign read_17d[19] = data_0n[19];
  assign read_17d[20] = data_0n[20];
  assign read_17d[21] = data_0n[21];
  assign read_17d[22] = data_0n[22];
  assign read_17d[23] = data_0n[23];
  assign read_17d[24] = data_0n[24];
  assign read_17d[25] = data_0n[25];
  assign read_17d[26] = data_0n[26];
  assign read_17d[27] = data_0n[27];
  assign read_17d[28] = data_0n[28];
  assign read_17d[29] = data_0n[29];
  assign read_17d[30] = data_0n[30];
  assign read_17d[31] = data_0n[31];
  assign read_17d[32] = data_0n[32];
  assign read_16d[0] = data_0n[0];
  assign read_16d[1] = data_0n[1];
  assign read_16d[2] = data_0n[2];
  assign read_16d[3] = data_0n[3];
  assign read_16d[4] = data_0n[4];
  assign read_16d[5] = data_0n[5];
  assign read_16d[6] = data_0n[6];
  assign read_16d[7] = data_0n[7];
  assign read_16d[8] = data_0n[8];
  assign read_16d[9] = data_0n[9];
  assign read_16d[10] = data_0n[10];
  assign read_16d[11] = data_0n[11];
  assign read_16d[12] = data_0n[12];
  assign read_16d[13] = data_0n[13];
  assign read_16d[14] = data_0n[14];
  assign read_16d[15] = data_0n[15];
  assign read_16d[16] = data_0n[16];
  assign read_16d[17] = data_0n[17];
  assign read_16d[18] = data_0n[18];
  assign read_16d[19] = data_0n[19];
  assign read_16d[20] = data_0n[20];
  assign read_16d[21] = data_0n[21];
  assign read_16d[22] = data_0n[22];
  assign read_16d[23] = data_0n[23];
  assign read_16d[24] = data_0n[24];
  assign read_16d[25] = data_0n[25];
  assign read_16d[26] = data_0n[26];
  assign read_16d[27] = data_0n[27];
  assign read_16d[28] = data_0n[28];
  assign read_16d[29] = data_0n[29];
  assign read_16d[30] = data_0n[30];
  assign read_16d[31] = data_0n[31];
  assign read_16d[32] = data_0n[32];
  assign read_15d[0] = data_0n[0];
  assign read_15d[1] = data_0n[1];
  assign read_15d[2] = data_0n[2];
  assign read_15d[3] = data_0n[3];
  assign read_15d[4] = data_0n[4];
  assign read_15d[5] = data_0n[5];
  assign read_15d[6] = data_0n[6];
  assign read_15d[7] = data_0n[7];
  assign read_15d[8] = data_0n[8];
  assign read_15d[9] = data_0n[9];
  assign read_15d[10] = data_0n[10];
  assign read_15d[11] = data_0n[11];
  assign read_15d[12] = data_0n[12];
  assign read_15d[13] = data_0n[13];
  assign read_15d[14] = data_0n[14];
  assign read_15d[15] = data_0n[15];
  assign read_15d[16] = data_0n[16];
  assign read_15d[17] = data_0n[17];
  assign read_15d[18] = data_0n[18];
  assign read_15d[19] = data_0n[19];
  assign read_15d[20] = data_0n[20];
  assign read_15d[21] = data_0n[21];
  assign read_15d[22] = data_0n[22];
  assign read_15d[23] = data_0n[23];
  assign read_15d[24] = data_0n[24];
  assign read_15d[25] = data_0n[25];
  assign read_15d[26] = data_0n[26];
  assign read_15d[27] = data_0n[27];
  assign read_15d[28] = data_0n[28];
  assign read_15d[29] = data_0n[29];
  assign read_15d[30] = data_0n[30];
  assign read_15d[31] = data_0n[31];
  assign read_15d[32] = data_0n[32];
  assign read_14d[0] = data_0n[0];
  assign read_14d[1] = data_0n[1];
  assign read_14d[2] = data_0n[2];
  assign read_14d[3] = data_0n[3];
  assign read_14d[4] = data_0n[4];
  assign read_14d[5] = data_0n[5];
  assign read_14d[6] = data_0n[6];
  assign read_14d[7] = data_0n[7];
  assign read_14d[8] = data_0n[8];
  assign read_14d[9] = data_0n[9];
  assign read_14d[10] = data_0n[10];
  assign read_14d[11] = data_0n[11];
  assign read_14d[12] = data_0n[12];
  assign read_14d[13] = data_0n[13];
  assign read_14d[14] = data_0n[14];
  assign read_14d[15] = data_0n[15];
  assign read_14d[16] = data_0n[16];
  assign read_14d[17] = data_0n[17];
  assign read_14d[18] = data_0n[18];
  assign read_14d[19] = data_0n[19];
  assign read_14d[20] = data_0n[20];
  assign read_14d[21] = data_0n[21];
  assign read_14d[22] = data_0n[22];
  assign read_14d[23] = data_0n[23];
  assign read_14d[24] = data_0n[24];
  assign read_14d[25] = data_0n[25];
  assign read_14d[26] = data_0n[26];
  assign read_14d[27] = data_0n[27];
  assign read_14d[28] = data_0n[28];
  assign read_14d[29] = data_0n[29];
  assign read_14d[30] = data_0n[30];
  assign read_14d[31] = data_0n[31];
  assign read_14d[32] = data_0n[32];
  assign read_13d = data_0n[0];
  assign read_12d = data_0n[1];
  assign read_11d = data_0n[0];
  assign read_10d = data_0n[1];
  assign read_9d = data_0n[32];
  assign read_8d[0] = data_0n[1];
  assign read_8d[1] = data_0n[2];
  assign read_8d[2] = data_0n[3];
  assign read_8d[3] = data_0n[4];
  assign read_8d[4] = data_0n[5];
  assign read_8d[5] = data_0n[6];
  assign read_8d[6] = data_0n[7];
  assign read_8d[7] = data_0n[8];
  assign read_8d[8] = data_0n[9];
  assign read_8d[9] = data_0n[10];
  assign read_8d[10] = data_0n[11];
  assign read_8d[11] = data_0n[12];
  assign read_8d[12] = data_0n[13];
  assign read_8d[13] = data_0n[14];
  assign read_8d[14] = data_0n[15];
  assign read_8d[15] = data_0n[16];
  assign read_8d[16] = data_0n[17];
  assign read_8d[17] = data_0n[18];
  assign read_8d[18] = data_0n[19];
  assign read_8d[19] = data_0n[20];
  assign read_8d[20] = data_0n[21];
  assign read_8d[21] = data_0n[22];
  assign read_8d[22] = data_0n[23];
  assign read_8d[23] = data_0n[24];
  assign read_8d[24] = data_0n[25];
  assign read_8d[25] = data_0n[26];
  assign read_8d[26] = data_0n[27];
  assign read_8d[27] = data_0n[28];
  assign read_8d[28] = data_0n[29];
  assign read_8d[29] = data_0n[30];
  assign read_8d[30] = data_0n[31];
  assign read_8d[31] = data_0n[32];
  assign read_7d[0] = data_0n[0];
  assign read_7d[1] = data_0n[1];
  assign read_7d[2] = data_0n[2];
  assign read_7d[3] = data_0n[3];
  assign read_7d[4] = data_0n[4];
  assign read_7d[5] = data_0n[5];
  assign read_7d[6] = data_0n[6];
  assign read_7d[7] = data_0n[7];
  assign read_7d[8] = data_0n[8];
  assign read_7d[9] = data_0n[9];
  assign read_7d[10] = data_0n[10];
  assign read_7d[11] = data_0n[11];
  assign read_7d[12] = data_0n[12];
  assign read_7d[13] = data_0n[13];
  assign read_7d[14] = data_0n[14];
  assign read_7d[15] = data_0n[15];
  assign read_7d[16] = data_0n[16];
  assign read_7d[17] = data_0n[17];
  assign read_7d[18] = data_0n[18];
  assign read_7d[19] = data_0n[19];
  assign read_7d[20] = data_0n[20];
  assign read_7d[21] = data_0n[21];
  assign read_7d[22] = data_0n[22];
  assign read_7d[23] = data_0n[23];
  assign read_7d[24] = data_0n[24];
  assign read_7d[25] = data_0n[25];
  assign read_7d[26] = data_0n[26];
  assign read_7d[27] = data_0n[27];
  assign read_7d[28] = data_0n[28];
  assign read_7d[29] = data_0n[29];
  assign read_7d[30] = data_0n[30];
  assign read_7d[31] = data_0n[31];
  assign read_7d[32] = data_0n[32];
  assign read_6d[0] = data_0n[0];
  assign read_6d[1] = data_0n[1];
  assign read_6d[2] = data_0n[2];
  assign read_6d[3] = data_0n[3];
  assign read_6d[4] = data_0n[4];
  assign read_6d[5] = data_0n[5];
  assign read_6d[6] = data_0n[6];
  assign read_6d[7] = data_0n[7];
  assign read_6d[8] = data_0n[8];
  assign read_6d[9] = data_0n[9];
  assign read_6d[10] = data_0n[10];
  assign read_6d[11] = data_0n[11];
  assign read_6d[12] = data_0n[12];
  assign read_6d[13] = data_0n[13];
  assign read_6d[14] = data_0n[14];
  assign read_6d[15] = data_0n[15];
  assign read_6d[16] = data_0n[16];
  assign read_6d[17] = data_0n[17];
  assign read_6d[18] = data_0n[18];
  assign read_6d[19] = data_0n[19];
  assign read_6d[20] = data_0n[20];
  assign read_6d[21] = data_0n[21];
  assign read_6d[22] = data_0n[22];
  assign read_6d[23] = data_0n[23];
  assign read_6d[24] = data_0n[24];
  assign read_6d[25] = data_0n[25];
  assign read_6d[26] = data_0n[26];
  assign read_6d[27] = data_0n[27];
  assign read_6d[28] = data_0n[28];
  assign read_6d[29] = data_0n[29];
  assign read_6d[30] = data_0n[30];
  assign read_6d[31] = data_0n[31];
  assign read_6d[32] = data_0n[32];
  assign read_5d[0] = data_0n[0];
  assign read_5d[1] = data_0n[1];
  assign read_5d[2] = data_0n[2];
  assign read_5d[3] = data_0n[3];
  assign read_5d[4] = data_0n[4];
  assign read_5d[5] = data_0n[5];
  assign read_5d[6] = data_0n[6];
  assign read_5d[7] = data_0n[7];
  assign read_5d[8] = data_0n[8];
  assign read_5d[9] = data_0n[9];
  assign read_5d[10] = data_0n[10];
  assign read_5d[11] = data_0n[11];
  assign read_5d[12] = data_0n[12];
  assign read_5d[13] = data_0n[13];
  assign read_5d[14] = data_0n[14];
  assign read_5d[15] = data_0n[15];
  assign read_5d[16] = data_0n[16];
  assign read_5d[17] = data_0n[17];
  assign read_5d[18] = data_0n[18];
  assign read_5d[19] = data_0n[19];
  assign read_5d[20] = data_0n[20];
  assign read_5d[21] = data_0n[21];
  assign read_5d[22] = data_0n[22];
  assign read_5d[23] = data_0n[23];
  assign read_5d[24] = data_0n[24];
  assign read_5d[25] = data_0n[25];
  assign read_5d[26] = data_0n[26];
  assign read_5d[27] = data_0n[27];
  assign read_5d[28] = data_0n[28];
  assign read_5d[29] = data_0n[29];
  assign read_5d[30] = data_0n[30];
  assign read_5d[31] = data_0n[31];
  assign read_5d[32] = data_0n[32];
  assign read_4d[0] = data_0n[0];
  assign read_4d[1] = data_0n[1];
  assign read_4d[2] = data_0n[2];
  assign read_4d[3] = data_0n[3];
  assign read_4d[4] = data_0n[4];
  assign read_4d[5] = data_0n[5];
  assign read_4d[6] = data_0n[6];
  assign read_4d[7] = data_0n[7];
  assign read_4d[8] = data_0n[8];
  assign read_4d[9] = data_0n[9];
  assign read_4d[10] = data_0n[10];
  assign read_4d[11] = data_0n[11];
  assign read_4d[12] = data_0n[12];
  assign read_4d[13] = data_0n[13];
  assign read_4d[14] = data_0n[14];
  assign read_4d[15] = data_0n[15];
  assign read_4d[16] = data_0n[16];
  assign read_4d[17] = data_0n[17];
  assign read_4d[18] = data_0n[18];
  assign read_4d[19] = data_0n[19];
  assign read_4d[20] = data_0n[20];
  assign read_4d[21] = data_0n[21];
  assign read_4d[22] = data_0n[22];
  assign read_4d[23] = data_0n[23];
  assign read_4d[24] = data_0n[24];
  assign read_4d[25] = data_0n[25];
  assign read_4d[26] = data_0n[26];
  assign read_4d[27] = data_0n[27];
  assign read_4d[28] = data_0n[28];
  assign read_4d[29] = data_0n[29];
  assign read_4d[30] = data_0n[30];
  assign read_4d[31] = data_0n[31];
  assign read_4d[32] = data_0n[32];
  assign read_3d = data_0n[0];
  assign read_2d = data_0n[1];
  assign read_1d = data_0n[0];
  assign read_0d = data_0n[1];
  LD1 I2897 (write_0d[0], bWriteReq_0n, data_0n[0]);
  LD1 I2898 (write_0d[1], bWriteReq_0n, data_0n[1]);
  LD1 I2899 (write_0d[2], bWriteReq_0n, data_0n[2]);
  LD1 I2900 (write_0d[3], bWriteReq_0n, data_0n[3]);
  LD1 I2901 (write_0d[4], bWriteReq_0n, data_0n[4]);
  LD1 I2902 (write_0d[5], bWriteReq_0n, data_0n[5]);
  LD1 I2903 (write_0d[6], bWriteReq_0n, data_0n[6]);
  LD1 I2904 (write_0d[7], bWriteReq_0n, data_0n[7]);
  LD1 I2905 (write_0d[8], bWriteReq_0n, data_0n[8]);
  LD1 I2906 (write_0d[9], bWriteReq_0n, data_0n[9]);
  LD1 I2907 (write_0d[10], bWriteReq_0n, data_0n[10]);
  LD1 I2908 (write_0d[11], bWriteReq_0n, data_0n[11]);
  LD1 I2909 (write_0d[12], bWriteReq_0n, data_0n[12]);
  LD1 I2910 (write_0d[13], bWriteReq_0n, data_0n[13]);
  LD1 I2911 (write_0d[14], bWriteReq_0n, data_0n[14]);
  LD1 I2912 (write_0d[15], bWriteReq_0n, data_0n[15]);
  LD1 I2913 (write_0d[16], bWriteReq_0n, data_0n[16]);
  LD1 I2914 (write_0d[17], bWriteReq_0n, data_0n[17]);
  LD1 I2915 (write_0d[18], bWriteReq_0n, data_0n[18]);
  LD1 I2916 (write_0d[19], bWriteReq_0n, data_0n[19]);
  LD1 I2917 (write_0d[20], bWriteReq_0n, data_0n[20]);
  LD1 I2918 (write_0d[21], bWriteReq_0n, data_0n[21]);
  LD1 I2919 (write_0d[22], bWriteReq_0n, data_0n[22]);
  LD1 I2920 (write_0d[23], bWriteReq_0n, data_0n[23]);
  LD1 I2921 (write_0d[24], bWriteReq_0n, data_0n[24]);
  LD1 I2922 (write_0d[25], bWriteReq_0n, data_0n[25]);
  LD1 I2923 (write_0d[26], bWriteReq_0n, data_0n[26]);
  LD1 I2924 (write_0d[27], bWriteReq_0n, data_0n[27]);
  LD1 I2925 (write_0d[28], bWriteReq_0n, data_0n[28]);
  LD1 I2926 (write_0d[29], bWriteReq_0n, data_0n[29]);
  LD1 I2927 (write_0d[30], bWriteReq_0n, data_0n[30]);
  LD1 I2928 (write_0d[31], bWriteReq_0n, data_0n[31]);
  LD1 I2929 (write_0d[32], bWriteReq_0n, data_0n[32]);
  IV I2930 (write_0a, nbWriteReq_0n);
  IV I2931 (nbWriteReq_0n, bWriteReq_0n);
  IV I2932 (bWriteReq_0n, nWriteReq_0n);
  IV I2933 (nWriteReq_0n, write_0r);
endmodule

module Balsa_booth__mul16 (
  activate_0r, activate_0a,
  x_0r, x_0a, x_0d,
  y_0r, y_0a, y_0d,
  z_0r, z_0a, z_0d
);
  input activate_0r;
  output activate_0a;
  output x_0r;
  input x_0a;
  input [15:0] x_0d;
  output y_0r;
  input y_0a;
  input [15:0] y_0d;
  output z_0r;
  input z_0a;
  output [31:0] z_0d;
  wire c895_r;
  wire c895_a;
  wire [32:0] c895_d;
  wire c894_r;
  wire c894_a;
  wire c893_r;
  wire c893_a;
  wire c892_r;
  wire c892_a;
  wire c891_r;
  wire c891_a;
  wire [15:0] c891_d;
  wire c890_r;
  wire c890_a;
  wire c889_r;
  wire c889_a;
  wire [15:0] c889_d;
  wire c888_r;
  wire c888_a;
  wire c887_r;
  wire c887_a;
  wire c886_r;
  wire c886_a;
  wire [32:0] c886_d;
  wire c885_r;
  wire c885_a;
  wire [32:0] c885_d;
  wire c884_r;
  wire c884_a;
  wire [16:0] c884_d;
  wire c883_r;
  wire c883_a;
  wire [15:0] c883_d;
  wire c882_r;
  wire c882_a;
  wire c881_r;
  wire c881_a;
  wire [32:0] c881_d;
  wire c880_r;
  wire c880_a;
  wire [32:0] c880_d;
  wire c879_r;
  wire c879_a;
  wire [16:0] c879_d;
  wire c878_r;
  wire c878_a;
  wire [15:0] c878_d;
  wire c877_r;
  wire c877_a;
  wire [15:0] c877_d;
  wire c876_r;
  wire c876_a;
  wire c875_r;
  wire c875_a;
  wire [32:0] c875_d;
  wire c874_r;
  wire c874_a;
  wire [32:0] c874_d;
  wire c873_r;
  wire c873_a;
  wire [16:0] c873_d;
  wire c872_r;
  wire c872_a;
  wire c872_d;
  wire c871_r;
  wire c871_a;
  wire [15:0] c871_d;
  wire c870_r;
  wire c870_a;
  wire c870_d;
  wire c869_r;
  wire c869_a;
  wire c869_d;
  wire c868_r;
  wire c868_a;
  wire c867_r;
  wire c867_a;
  wire c866_r;
  wire c866_a;
  wire c866_d;
  wire c865_r;
  wire c865_a;
  wire c864_r;
  wire c864_a;
  wire c864_d;
  wire c863_r;
  wire c863_a;
  wire c863_d;
  wire c862_r;
  wire c862_a;
  wire c862_d;
  wire c861_r;
  wire c861_a;
  wire c861_d;
  wire c860_r;
  wire c860_a;
  wire c860_d;
  wire c859_r;
  wire c859_a;
  wire [32:0] c859_d;
  wire c858_r;
  wire c858_a;
  wire [32:0] c858_d;
  wire c857_r;
  wire c857_a;
  wire c856_r;
  wire c856_a;
  wire c855_r;
  wire c855_a;
  wire c854_r;
  wire c854_a;
  wire [32:0] c854_d;
  wire c853_r;
  wire c853_a;
  wire [32:0] c853_d;
  wire c852_r;
  wire c852_a;
  wire [31:0] c852_d;
  wire c851_r;
  wire c851_a;
  wire [33:0] c851_d;
  wire c850_r;
  wire c850_a;
  wire [32:0] c850_d;
  wire c849_r;
  wire c849_a;
  wire [32:0] c849_d;
  wire c848_r;
  wire c848_a;
  wire c848_d;
  wire c847_r;
  wire c847_a;
  wire [33:0] c847_d;
  wire c846_r;
  wire c846_a;
  wire [32:0] c846_d;
  wire c845_r;
  wire c845_a;
  wire [32:0] c845_d;
  wire c844_r;
  wire c844_a;
  wire c844_d;
  wire c843_r;
  wire c843_a;
  wire c843_d;
  wire c842_r;
  wire c842_a;
  wire c842_d;
  wire c841_r;
  wire c841_a;
  wire c841_d;
  wire c840_r;
  wire c840_a;
  wire [32:0] c840_d;
  wire c839_r;
  wire c839_a;
  wire [32:0] c839_d;
  wire c838_r;
  wire c838_a;
  wire c837_r;
  wire c837_a;
  wire c836_r;
  wire c836_a;
  wire c835_r;
  wire c835_a;
  wire [32:0] c835_d;
  wire c834_r;
  wire c834_a;
  wire [32:0] c834_d;
  wire c833_r;
  wire c833_a;
  wire [31:0] c833_d;
  wire c832_r;
  wire c832_a;
  wire [33:0] c832_d;
  wire c831_r;
  wire c831_a;
  wire [32:0] c831_d;
  wire c830_r;
  wire c830_a;
  wire [32:0] c830_d;
  wire c829_r;
  wire c829_a;
  wire c829_d;
  wire c828_r;
  wire c828_a;
  wire [33:0] c828_d;
  wire c827_r;
  wire c827_a;
  wire [32:0] c827_d;
  wire c826_r;
  wire c826_a;
  wire [32:0] c826_d;
  wire c825_r;
  wire c825_a;
  wire [32:0] c825_d;
  wire c824_r;
  wire c824_a;
  wire [32:0] c824_d;
  wire c823_r;
  wire c823_a;
  wire c822_r;
  wire c822_a;
  wire c821_r;
  wire c821_a;
  wire c820_r;
  wire c820_a;
  wire [32:0] c820_d;
  wire c819_r;
  wire c819_a;
  wire [32:0] c819_d;
  wire c818_r;
  wire c818_a;
  wire [31:0] c818_d;
  wire c817_r;
  wire c817_a;
  wire c817_d;
  wire c816_r;
  wire c816_a;
  wire c816_d;
  wire c815_r;
  wire c815_a;
  wire c815_d;
  wire c814_r;
  wire c814_a;
  wire c813_r;
  wire c813_a;
  wire c812_r;
  wire c812_a;
  wire c812_d;
  wire c811_r;
  wire c811_a;
  wire c810_r;
  wire c810_a;
  wire c810_d;
  wire c809_r;
  wire c809_a;
  wire c809_d;
  wire c808_r;
  wire c808_a;
  wire c808_d;
  wire c807_r;
  wire c807_a;
  wire c807_d;
  wire c806_r;
  wire c806_a;
  wire c806_d;
  wire c805_r;
  wire c805_a;
  wire [32:0] c805_d;
  wire c804_r;
  wire c804_a;
  wire [32:0] c804_d;
  wire c803_r;
  wire c803_a;
  wire c802_r;
  wire c802_a;
  wire c801_r;
  wire c801_a;
  wire c800_r;
  wire c800_a;
  wire [32:0] c800_d;
  wire c799_r;
  wire c799_a;
  wire [32:0] c799_d;
  wire c798_r;
  wire c798_a;
  wire [31:0] c798_d;
  wire c797_r;
  wire c797_a;
  wire [33:0] c797_d;
  wire c796_r;
  wire c796_a;
  wire [32:0] c796_d;
  wire c795_r;
  wire c795_a;
  wire [32:0] c795_d;
  wire c794_r;
  wire c794_a;
  wire c794_d;
  wire c793_r;
  wire c793_a;
  wire [33:0] c793_d;
  wire c792_r;
  wire c792_a;
  wire [32:0] c792_d;
  wire c791_r;
  wire c791_a;
  wire [32:0] c791_d;
  wire c790_r;
  wire c790_a;
  wire c790_d;
  wire c789_r;
  wire c789_a;
  wire c789_d;
  wire c788_r;
  wire c788_a;
  wire c788_d;
  wire c787_r;
  wire c787_a;
  wire c787_d;
  wire c786_r;
  wire c786_a;
  wire [32:0] c786_d;
  wire c785_r;
  wire c785_a;
  wire [32:0] c785_d;
  wire c784_r;
  wire c784_a;
  wire c783_r;
  wire c783_a;
  wire c782_r;
  wire c782_a;
  wire c781_r;
  wire c781_a;
  wire [32:0] c781_d;
  wire c780_r;
  wire c780_a;
  wire [32:0] c780_d;
  wire c779_r;
  wire c779_a;
  wire [31:0] c779_d;
  wire c778_r;
  wire c778_a;
  wire [33:0] c778_d;
  wire c777_r;
  wire c777_a;
  wire [32:0] c777_d;
  wire c776_r;
  wire c776_a;
  wire [32:0] c776_d;
  wire c775_r;
  wire c775_a;
  wire c775_d;
  wire c774_r;
  wire c774_a;
  wire [33:0] c774_d;
  wire c773_r;
  wire c773_a;
  wire [32:0] c773_d;
  wire c772_r;
  wire c772_a;
  wire [32:0] c772_d;
  wire c771_r;
  wire c771_a;
  wire [32:0] c771_d;
  wire c770_r;
  wire c770_a;
  wire [32:0] c770_d;
  wire c769_r;
  wire c769_a;
  wire c768_r;
  wire c768_a;
  wire c767_r;
  wire c767_a;
  wire c766_r;
  wire c766_a;
  wire [32:0] c766_d;
  wire c765_r;
  wire c765_a;
  wire [32:0] c765_d;
  wire c764_r;
  wire c764_a;
  wire [31:0] c764_d;
  wire c763_r;
  wire c763_a;
  wire c763_d;
  wire c762_r;
  wire c762_a;
  wire c762_d;
  wire c761_r;
  wire c761_a;
  wire c761_d;
  wire c760_r;
  wire c760_a;
  wire c759_r;
  wire c759_a;
  wire c758_r;
  wire c758_a;
  wire c758_d;
  wire c757_r;
  wire c757_a;
  wire c756_r;
  wire c756_a;
  wire c756_d;
  wire c755_r;
  wire c755_a;
  wire c755_d;
  wire c754_r;
  wire c754_a;
  wire c754_d;
  wire c753_r;
  wire c753_a;
  wire c753_d;
  wire c752_r;
  wire c752_a;
  wire c752_d;
  wire c751_r;
  wire c751_a;
  wire [32:0] c751_d;
  wire c750_r;
  wire c750_a;
  wire [32:0] c750_d;
  wire c749_r;
  wire c749_a;
  wire c748_r;
  wire c748_a;
  wire c747_r;
  wire c747_a;
  wire c746_r;
  wire c746_a;
  wire [32:0] c746_d;
  wire c745_r;
  wire c745_a;
  wire [32:0] c745_d;
  wire c744_r;
  wire c744_a;
  wire [31:0] c744_d;
  wire c743_r;
  wire c743_a;
  wire [33:0] c743_d;
  wire c742_r;
  wire c742_a;
  wire [32:0] c742_d;
  wire c741_r;
  wire c741_a;
  wire [32:0] c741_d;
  wire c740_r;
  wire c740_a;
  wire c740_d;
  wire c739_r;
  wire c739_a;
  wire [33:0] c739_d;
  wire c738_r;
  wire c738_a;
  wire [32:0] c738_d;
  wire c737_r;
  wire c737_a;
  wire [32:0] c737_d;
  wire c736_r;
  wire c736_a;
  wire c736_d;
  wire c735_r;
  wire c735_a;
  wire c735_d;
  wire c734_r;
  wire c734_a;
  wire c734_d;
  wire c733_r;
  wire c733_a;
  wire c733_d;
  wire c732_r;
  wire c732_a;
  wire [32:0] c732_d;
  wire c731_r;
  wire c731_a;
  wire [32:0] c731_d;
  wire c730_r;
  wire c730_a;
  wire c729_r;
  wire c729_a;
  wire c728_r;
  wire c728_a;
  wire c727_r;
  wire c727_a;
  wire [32:0] c727_d;
  wire c726_r;
  wire c726_a;
  wire [32:0] c726_d;
  wire c725_r;
  wire c725_a;
  wire [31:0] c725_d;
  wire c724_r;
  wire c724_a;
  wire [33:0] c724_d;
  wire c723_r;
  wire c723_a;
  wire [32:0] c723_d;
  wire c722_r;
  wire c722_a;
  wire [32:0] c722_d;
  wire c721_r;
  wire c721_a;
  wire c721_d;
  wire c720_r;
  wire c720_a;
  wire [33:0] c720_d;
  wire c719_r;
  wire c719_a;
  wire [32:0] c719_d;
  wire c718_r;
  wire c718_a;
  wire [32:0] c718_d;
  wire c717_r;
  wire c717_a;
  wire [32:0] c717_d;
  wire c716_r;
  wire c716_a;
  wire [32:0] c716_d;
  wire c715_r;
  wire c715_a;
  wire c714_r;
  wire c714_a;
  wire c713_r;
  wire c713_a;
  wire c712_r;
  wire c712_a;
  wire [32:0] c712_d;
  wire c711_r;
  wire c711_a;
  wire [32:0] c711_d;
  wire c710_r;
  wire c710_a;
  wire [31:0] c710_d;
  wire c709_r;
  wire c709_a;
  wire c709_d;
  wire c708_r;
  wire c708_a;
  wire c708_d;
  wire c707_r;
  wire c707_a;
  wire c707_d;
  wire c706_r;
  wire c706_a;
  wire c705_r;
  wire c705_a;
  wire c704_r;
  wire c704_a;
  wire c704_d;
  wire c703_r;
  wire c703_a;
  wire c702_r;
  wire c702_a;
  wire c702_d;
  wire c701_r;
  wire c701_a;
  wire c701_d;
  wire c700_r;
  wire c700_a;
  wire c700_d;
  wire c699_r;
  wire c699_a;
  wire c699_d;
  wire c698_r;
  wire c698_a;
  wire c698_d;
  wire c697_r;
  wire c697_a;
  wire [32:0] c697_d;
  wire c696_r;
  wire c696_a;
  wire [32:0] c696_d;
  wire c695_r;
  wire c695_a;
  wire c694_r;
  wire c694_a;
  wire c693_r;
  wire c693_a;
  wire c692_r;
  wire c692_a;
  wire [32:0] c692_d;
  wire c691_r;
  wire c691_a;
  wire [32:0] c691_d;
  wire c690_r;
  wire c690_a;
  wire [31:0] c690_d;
  wire c689_r;
  wire c689_a;
  wire [33:0] c689_d;
  wire c688_r;
  wire c688_a;
  wire [32:0] c688_d;
  wire c687_r;
  wire c687_a;
  wire [32:0] c687_d;
  wire c686_r;
  wire c686_a;
  wire c686_d;
  wire c685_r;
  wire c685_a;
  wire [33:0] c685_d;
  wire c684_r;
  wire c684_a;
  wire [32:0] c684_d;
  wire c683_r;
  wire c683_a;
  wire [32:0] c683_d;
  wire c682_r;
  wire c682_a;
  wire c682_d;
  wire c681_r;
  wire c681_a;
  wire c681_d;
  wire c680_r;
  wire c680_a;
  wire c680_d;
  wire c679_r;
  wire c679_a;
  wire c679_d;
  wire c678_r;
  wire c678_a;
  wire [32:0] c678_d;
  wire c677_r;
  wire c677_a;
  wire [32:0] c677_d;
  wire c676_r;
  wire c676_a;
  wire c675_r;
  wire c675_a;
  wire c674_r;
  wire c674_a;
  wire c673_r;
  wire c673_a;
  wire [32:0] c673_d;
  wire c672_r;
  wire c672_a;
  wire [32:0] c672_d;
  wire c671_r;
  wire c671_a;
  wire [31:0] c671_d;
  wire c670_r;
  wire c670_a;
  wire [33:0] c670_d;
  wire c669_r;
  wire c669_a;
  wire [32:0] c669_d;
  wire c668_r;
  wire c668_a;
  wire [32:0] c668_d;
  wire c667_r;
  wire c667_a;
  wire c667_d;
  wire c666_r;
  wire c666_a;
  wire [33:0] c666_d;
  wire c665_r;
  wire c665_a;
  wire [32:0] c665_d;
  wire c664_r;
  wire c664_a;
  wire [32:0] c664_d;
  wire c663_r;
  wire c663_a;
  wire [32:0] c663_d;
  wire c662_r;
  wire c662_a;
  wire [32:0] c662_d;
  wire c661_r;
  wire c661_a;
  wire c660_r;
  wire c660_a;
  wire c659_r;
  wire c659_a;
  wire c658_r;
  wire c658_a;
  wire [32:0] c658_d;
  wire c657_r;
  wire c657_a;
  wire [32:0] c657_d;
  wire c656_r;
  wire c656_a;
  wire [31:0] c656_d;
  wire c655_r;
  wire c655_a;
  wire c655_d;
  wire c654_r;
  wire c654_a;
  wire c654_d;
  wire c653_r;
  wire c653_a;
  wire c653_d;
  wire c652_r;
  wire c652_a;
  wire c651_r;
  wire c651_a;
  wire c650_r;
  wire c650_a;
  wire c650_d;
  wire c649_r;
  wire c649_a;
  wire c648_r;
  wire c648_a;
  wire c648_d;
  wire c647_r;
  wire c647_a;
  wire c647_d;
  wire c646_r;
  wire c646_a;
  wire c646_d;
  wire c645_r;
  wire c645_a;
  wire c645_d;
  wire c644_r;
  wire c644_a;
  wire c644_d;
  wire c643_r;
  wire c643_a;
  wire [32:0] c643_d;
  wire c642_r;
  wire c642_a;
  wire [32:0] c642_d;
  wire c641_r;
  wire c641_a;
  wire c640_r;
  wire c640_a;
  wire c639_r;
  wire c639_a;
  wire c638_r;
  wire c638_a;
  wire [32:0] c638_d;
  wire c637_r;
  wire c637_a;
  wire [32:0] c637_d;
  wire c636_r;
  wire c636_a;
  wire [31:0] c636_d;
  wire c635_r;
  wire c635_a;
  wire [33:0] c635_d;
  wire c634_r;
  wire c634_a;
  wire [32:0] c634_d;
  wire c633_r;
  wire c633_a;
  wire [32:0] c633_d;
  wire c632_r;
  wire c632_a;
  wire c632_d;
  wire c631_r;
  wire c631_a;
  wire [33:0] c631_d;
  wire c630_r;
  wire c630_a;
  wire [32:0] c630_d;
  wire c629_r;
  wire c629_a;
  wire [32:0] c629_d;
  wire c628_r;
  wire c628_a;
  wire c628_d;
  wire c627_r;
  wire c627_a;
  wire c627_d;
  wire c626_r;
  wire c626_a;
  wire c626_d;
  wire c625_r;
  wire c625_a;
  wire c625_d;
  wire c624_r;
  wire c624_a;
  wire [32:0] c624_d;
  wire c623_r;
  wire c623_a;
  wire [32:0] c623_d;
  wire c622_r;
  wire c622_a;
  wire c621_r;
  wire c621_a;
  wire c620_r;
  wire c620_a;
  wire c619_r;
  wire c619_a;
  wire [32:0] c619_d;
  wire c618_r;
  wire c618_a;
  wire [32:0] c618_d;
  wire c617_r;
  wire c617_a;
  wire [31:0] c617_d;
  wire c616_r;
  wire c616_a;
  wire [33:0] c616_d;
  wire c615_r;
  wire c615_a;
  wire [32:0] c615_d;
  wire c614_r;
  wire c614_a;
  wire [32:0] c614_d;
  wire c613_r;
  wire c613_a;
  wire c613_d;
  wire c612_r;
  wire c612_a;
  wire [33:0] c612_d;
  wire c611_r;
  wire c611_a;
  wire [32:0] c611_d;
  wire c610_r;
  wire c610_a;
  wire [32:0] c610_d;
  wire c609_r;
  wire c609_a;
  wire [32:0] c609_d;
  wire c608_r;
  wire c608_a;
  wire [32:0] c608_d;
  wire c607_r;
  wire c607_a;
  wire c606_r;
  wire c606_a;
  wire c605_r;
  wire c605_a;
  wire c604_r;
  wire c604_a;
  wire [32:0] c604_d;
  wire c603_r;
  wire c603_a;
  wire [32:0] c603_d;
  wire c602_r;
  wire c602_a;
  wire [31:0] c602_d;
  wire c601_r;
  wire c601_a;
  wire c601_d;
  wire c600_r;
  wire c600_a;
  wire c600_d;
  wire c599_r;
  wire c599_a;
  wire c599_d;
  wire c598_r;
  wire c598_a;
  wire c597_r;
  wire c597_a;
  wire c596_r;
  wire c596_a;
  wire c596_d;
  wire c595_r;
  wire c595_a;
  wire c594_r;
  wire c594_a;
  wire c594_d;
  wire c593_r;
  wire c593_a;
  wire c593_d;
  wire c592_r;
  wire c592_a;
  wire c592_d;
  wire c591_r;
  wire c591_a;
  wire c591_d;
  wire c590_r;
  wire c590_a;
  wire c590_d;
  wire c589_r;
  wire c589_a;
  wire [32:0] c589_d;
  wire c588_r;
  wire c588_a;
  wire [32:0] c588_d;
  wire c587_r;
  wire c587_a;
  wire c586_r;
  wire c586_a;
  wire c585_r;
  wire c585_a;
  wire c584_r;
  wire c584_a;
  wire [32:0] c584_d;
  wire c583_r;
  wire c583_a;
  wire [32:0] c583_d;
  wire c582_r;
  wire c582_a;
  wire [31:0] c582_d;
  wire c581_r;
  wire c581_a;
  wire [33:0] c581_d;
  wire c580_r;
  wire c580_a;
  wire [32:0] c580_d;
  wire c579_r;
  wire c579_a;
  wire [32:0] c579_d;
  wire c578_r;
  wire c578_a;
  wire c578_d;
  wire c577_r;
  wire c577_a;
  wire [33:0] c577_d;
  wire c576_r;
  wire c576_a;
  wire [32:0] c576_d;
  wire c575_r;
  wire c575_a;
  wire [32:0] c575_d;
  wire c574_r;
  wire c574_a;
  wire c574_d;
  wire c573_r;
  wire c573_a;
  wire c573_d;
  wire c572_r;
  wire c572_a;
  wire c572_d;
  wire c571_r;
  wire c571_a;
  wire c571_d;
  wire c570_r;
  wire c570_a;
  wire [32:0] c570_d;
  wire c569_r;
  wire c569_a;
  wire [32:0] c569_d;
  wire c568_r;
  wire c568_a;
  wire c567_r;
  wire c567_a;
  wire c566_r;
  wire c566_a;
  wire c565_r;
  wire c565_a;
  wire [32:0] c565_d;
  wire c564_r;
  wire c564_a;
  wire [32:0] c564_d;
  wire c563_r;
  wire c563_a;
  wire [31:0] c563_d;
  wire c562_r;
  wire c562_a;
  wire [33:0] c562_d;
  wire c561_r;
  wire c561_a;
  wire [32:0] c561_d;
  wire c560_r;
  wire c560_a;
  wire [32:0] c560_d;
  wire c559_r;
  wire c559_a;
  wire c559_d;
  wire c558_r;
  wire c558_a;
  wire [33:0] c558_d;
  wire c557_r;
  wire c557_a;
  wire [32:0] c557_d;
  wire c556_r;
  wire c556_a;
  wire [32:0] c556_d;
  wire c555_r;
  wire c555_a;
  wire [32:0] c555_d;
  wire c554_r;
  wire c554_a;
  wire [32:0] c554_d;
  wire c553_r;
  wire c553_a;
  wire c552_r;
  wire c552_a;
  wire c551_r;
  wire c551_a;
  wire c550_r;
  wire c550_a;
  wire [32:0] c550_d;
  wire c549_r;
  wire c549_a;
  wire [32:0] c549_d;
  wire c548_r;
  wire c548_a;
  wire [31:0] c548_d;
  wire c547_r;
  wire c547_a;
  wire c547_d;
  wire c546_r;
  wire c546_a;
  wire c546_d;
  wire c545_r;
  wire c545_a;
  wire c545_d;
  wire c544_r;
  wire c544_a;
  wire c543_r;
  wire c543_a;
  wire c542_r;
  wire c542_a;
  wire c542_d;
  wire c541_r;
  wire c541_a;
  wire c540_r;
  wire c540_a;
  wire c540_d;
  wire c539_r;
  wire c539_a;
  wire c539_d;
  wire c538_r;
  wire c538_a;
  wire c538_d;
  wire c537_r;
  wire c537_a;
  wire c537_d;
  wire c536_r;
  wire c536_a;
  wire c536_d;
  wire c535_r;
  wire c535_a;
  wire [32:0] c535_d;
  wire c534_r;
  wire c534_a;
  wire [32:0] c534_d;
  wire c533_r;
  wire c533_a;
  wire c532_r;
  wire c532_a;
  wire c531_r;
  wire c531_a;
  wire c530_r;
  wire c530_a;
  wire [32:0] c530_d;
  wire c529_r;
  wire c529_a;
  wire [32:0] c529_d;
  wire c528_r;
  wire c528_a;
  wire [31:0] c528_d;
  wire c527_r;
  wire c527_a;
  wire [33:0] c527_d;
  wire c526_r;
  wire c526_a;
  wire [32:0] c526_d;
  wire c525_r;
  wire c525_a;
  wire [32:0] c525_d;
  wire c524_r;
  wire c524_a;
  wire c524_d;
  wire c523_r;
  wire c523_a;
  wire [33:0] c523_d;
  wire c522_r;
  wire c522_a;
  wire [32:0] c522_d;
  wire c521_r;
  wire c521_a;
  wire [32:0] c521_d;
  wire c520_r;
  wire c520_a;
  wire c520_d;
  wire c519_r;
  wire c519_a;
  wire c519_d;
  wire c518_r;
  wire c518_a;
  wire c518_d;
  wire c517_r;
  wire c517_a;
  wire c517_d;
  wire c516_r;
  wire c516_a;
  wire [32:0] c516_d;
  wire c515_r;
  wire c515_a;
  wire [32:0] c515_d;
  wire c514_r;
  wire c514_a;
  wire c513_r;
  wire c513_a;
  wire c512_r;
  wire c512_a;
  wire c511_r;
  wire c511_a;
  wire [32:0] c511_d;
  wire c510_r;
  wire c510_a;
  wire [32:0] c510_d;
  wire c509_r;
  wire c509_a;
  wire [31:0] c509_d;
  wire c508_r;
  wire c508_a;
  wire [33:0] c508_d;
  wire c507_r;
  wire c507_a;
  wire [32:0] c507_d;
  wire c506_r;
  wire c506_a;
  wire [32:0] c506_d;
  wire c505_r;
  wire c505_a;
  wire c505_d;
  wire c504_r;
  wire c504_a;
  wire [33:0] c504_d;
  wire c503_r;
  wire c503_a;
  wire [32:0] c503_d;
  wire c502_r;
  wire c502_a;
  wire [32:0] c502_d;
  wire c501_r;
  wire c501_a;
  wire [32:0] c501_d;
  wire c500_r;
  wire c500_a;
  wire [32:0] c500_d;
  wire c499_r;
  wire c499_a;
  wire c498_r;
  wire c498_a;
  wire c497_r;
  wire c497_a;
  wire c496_r;
  wire c496_a;
  wire [32:0] c496_d;
  wire c495_r;
  wire c495_a;
  wire [32:0] c495_d;
  wire c494_r;
  wire c494_a;
  wire [31:0] c494_d;
  wire c493_r;
  wire c493_a;
  wire c493_d;
  wire c492_r;
  wire c492_a;
  wire c492_d;
  wire c491_r;
  wire c491_a;
  wire c491_d;
  wire c490_r;
  wire c490_a;
  wire c489_r;
  wire c489_a;
  wire c488_r;
  wire c488_a;
  wire c488_d;
  wire c487_r;
  wire c487_a;
  wire c486_r;
  wire c486_a;
  wire c486_d;
  wire c485_r;
  wire c485_a;
  wire c485_d;
  wire c484_r;
  wire c484_a;
  wire c484_d;
  wire c483_r;
  wire c483_a;
  wire c483_d;
  wire c482_r;
  wire c482_a;
  wire c482_d;
  wire c481_r;
  wire c481_a;
  wire [32:0] c481_d;
  wire c480_r;
  wire c480_a;
  wire [32:0] c480_d;
  wire c479_r;
  wire c479_a;
  wire c478_r;
  wire c478_a;
  wire c477_r;
  wire c477_a;
  wire c476_r;
  wire c476_a;
  wire [32:0] c476_d;
  wire c475_r;
  wire c475_a;
  wire [32:0] c475_d;
  wire c474_r;
  wire c474_a;
  wire [31:0] c474_d;
  wire c473_r;
  wire c473_a;
  wire [33:0] c473_d;
  wire c472_r;
  wire c472_a;
  wire [32:0] c472_d;
  wire c471_r;
  wire c471_a;
  wire [32:0] c471_d;
  wire c470_r;
  wire c470_a;
  wire c470_d;
  wire c469_r;
  wire c469_a;
  wire [33:0] c469_d;
  wire c468_r;
  wire c468_a;
  wire [32:0] c468_d;
  wire c467_r;
  wire c467_a;
  wire [32:0] c467_d;
  wire c466_r;
  wire c466_a;
  wire c466_d;
  wire c465_r;
  wire c465_a;
  wire c465_d;
  wire c464_r;
  wire c464_a;
  wire c464_d;
  wire c463_r;
  wire c463_a;
  wire c463_d;
  wire c462_r;
  wire c462_a;
  wire [32:0] c462_d;
  wire c461_r;
  wire c461_a;
  wire [32:0] c461_d;
  wire c460_r;
  wire c460_a;
  wire c459_r;
  wire c459_a;
  wire c458_r;
  wire c458_a;
  wire c457_r;
  wire c457_a;
  wire [32:0] c457_d;
  wire c456_r;
  wire c456_a;
  wire [32:0] c456_d;
  wire c455_r;
  wire c455_a;
  wire [31:0] c455_d;
  wire c454_r;
  wire c454_a;
  wire [33:0] c454_d;
  wire c453_r;
  wire c453_a;
  wire [32:0] c453_d;
  wire c452_r;
  wire c452_a;
  wire [32:0] c452_d;
  wire c451_r;
  wire c451_a;
  wire c451_d;
  wire c450_r;
  wire c450_a;
  wire [33:0] c450_d;
  wire c449_r;
  wire c449_a;
  wire [32:0] c449_d;
  wire c448_r;
  wire c448_a;
  wire [32:0] c448_d;
  wire c447_r;
  wire c447_a;
  wire [32:0] c447_d;
  wire c446_r;
  wire c446_a;
  wire [32:0] c446_d;
  wire c445_r;
  wire c445_a;
  wire c444_r;
  wire c444_a;
  wire c443_r;
  wire c443_a;
  wire c442_r;
  wire c442_a;
  wire [32:0] c442_d;
  wire c441_r;
  wire c441_a;
  wire [32:0] c441_d;
  wire c440_r;
  wire c440_a;
  wire [31:0] c440_d;
  wire c439_r;
  wire c439_a;
  wire c439_d;
  wire c438_r;
  wire c438_a;
  wire c438_d;
  wire c437_r;
  wire c437_a;
  wire c437_d;
  wire c436_r;
  wire c436_a;
  wire c435_r;
  wire c435_a;
  wire c434_r;
  wire c434_a;
  wire c434_d;
  wire c433_r;
  wire c433_a;
  wire c432_r;
  wire c432_a;
  wire c432_d;
  wire c431_r;
  wire c431_a;
  wire c431_d;
  wire c430_r;
  wire c430_a;
  wire c430_d;
  wire c429_r;
  wire c429_a;
  wire c429_d;
  wire c428_r;
  wire c428_a;
  wire c428_d;
  wire c427_r;
  wire c427_a;
  wire [32:0] c427_d;
  wire c426_r;
  wire c426_a;
  wire [32:0] c426_d;
  wire c425_r;
  wire c425_a;
  wire c424_r;
  wire c424_a;
  wire c423_r;
  wire c423_a;
  wire c422_r;
  wire c422_a;
  wire [32:0] c422_d;
  wire c421_r;
  wire c421_a;
  wire [32:0] c421_d;
  wire c420_r;
  wire c420_a;
  wire [31:0] c420_d;
  wire c419_r;
  wire c419_a;
  wire [33:0] c419_d;
  wire c418_r;
  wire c418_a;
  wire [32:0] c418_d;
  wire c417_r;
  wire c417_a;
  wire [32:0] c417_d;
  wire c416_r;
  wire c416_a;
  wire c416_d;
  wire c415_r;
  wire c415_a;
  wire [33:0] c415_d;
  wire c414_r;
  wire c414_a;
  wire [32:0] c414_d;
  wire c413_r;
  wire c413_a;
  wire [32:0] c413_d;
  wire c412_r;
  wire c412_a;
  wire c412_d;
  wire c411_r;
  wire c411_a;
  wire c411_d;
  wire c410_r;
  wire c410_a;
  wire c410_d;
  wire c409_r;
  wire c409_a;
  wire c409_d;
  wire c408_r;
  wire c408_a;
  wire [32:0] c408_d;
  wire c407_r;
  wire c407_a;
  wire [32:0] c407_d;
  wire c406_r;
  wire c406_a;
  wire c405_r;
  wire c405_a;
  wire c404_r;
  wire c404_a;
  wire c403_r;
  wire c403_a;
  wire [32:0] c403_d;
  wire c402_r;
  wire c402_a;
  wire [32:0] c402_d;
  wire c401_r;
  wire c401_a;
  wire [31:0] c401_d;
  wire c400_r;
  wire c400_a;
  wire [33:0] c400_d;
  wire c399_r;
  wire c399_a;
  wire [32:0] c399_d;
  wire c398_r;
  wire c398_a;
  wire [32:0] c398_d;
  wire c397_r;
  wire c397_a;
  wire c397_d;
  wire c396_r;
  wire c396_a;
  wire [33:0] c396_d;
  wire c395_r;
  wire c395_a;
  wire [32:0] c395_d;
  wire c394_r;
  wire c394_a;
  wire [32:0] c394_d;
  wire c393_r;
  wire c393_a;
  wire [32:0] c393_d;
  wire c392_r;
  wire c392_a;
  wire [32:0] c392_d;
  wire c391_r;
  wire c391_a;
  wire c390_r;
  wire c390_a;
  wire c389_r;
  wire c389_a;
  wire c388_r;
  wire c388_a;
  wire [32:0] c388_d;
  wire c387_r;
  wire c387_a;
  wire [32:0] c387_d;
  wire c386_r;
  wire c386_a;
  wire [31:0] c386_d;
  wire c385_r;
  wire c385_a;
  wire c385_d;
  wire c384_r;
  wire c384_a;
  wire c384_d;
  wire c383_r;
  wire c383_a;
  wire c383_d;
  wire c382_r;
  wire c382_a;
  wire c381_r;
  wire c381_a;
  wire c380_r;
  wire c380_a;
  wire c380_d;
  wire c379_r;
  wire c379_a;
  wire c378_r;
  wire c378_a;
  wire c378_d;
  wire c377_r;
  wire c377_a;
  wire c377_d;
  wire c376_r;
  wire c376_a;
  wire c376_d;
  wire c375_r;
  wire c375_a;
  wire c375_d;
  wire c374_r;
  wire c374_a;
  wire c374_d;
  wire c373_r;
  wire c373_a;
  wire [32:0] c373_d;
  wire c372_r;
  wire c372_a;
  wire [32:0] c372_d;
  wire c371_r;
  wire c371_a;
  wire c370_r;
  wire c370_a;
  wire c369_r;
  wire c369_a;
  wire c368_r;
  wire c368_a;
  wire [32:0] c368_d;
  wire c367_r;
  wire c367_a;
  wire [32:0] c367_d;
  wire c366_r;
  wire c366_a;
  wire [31:0] c366_d;
  wire c365_r;
  wire c365_a;
  wire [33:0] c365_d;
  wire c364_r;
  wire c364_a;
  wire [32:0] c364_d;
  wire c363_r;
  wire c363_a;
  wire [32:0] c363_d;
  wire c362_r;
  wire c362_a;
  wire c362_d;
  wire c361_r;
  wire c361_a;
  wire [33:0] c361_d;
  wire c360_r;
  wire c360_a;
  wire [32:0] c360_d;
  wire c359_r;
  wire c359_a;
  wire [32:0] c359_d;
  wire c358_r;
  wire c358_a;
  wire c358_d;
  wire c357_r;
  wire c357_a;
  wire c357_d;
  wire c356_r;
  wire c356_a;
  wire c356_d;
  wire c355_r;
  wire c355_a;
  wire c355_d;
  wire c354_r;
  wire c354_a;
  wire [32:0] c354_d;
  wire c353_r;
  wire c353_a;
  wire [32:0] c353_d;
  wire c352_r;
  wire c352_a;
  wire c351_r;
  wire c351_a;
  wire c350_r;
  wire c350_a;
  wire c349_r;
  wire c349_a;
  wire [32:0] c349_d;
  wire c348_r;
  wire c348_a;
  wire [32:0] c348_d;
  wire c347_r;
  wire c347_a;
  wire [31:0] c347_d;
  wire c346_r;
  wire c346_a;
  wire [33:0] c346_d;
  wire c345_r;
  wire c345_a;
  wire [32:0] c345_d;
  wire c344_r;
  wire c344_a;
  wire [32:0] c344_d;
  wire c343_r;
  wire c343_a;
  wire c343_d;
  wire c342_r;
  wire c342_a;
  wire [33:0] c342_d;
  wire c341_r;
  wire c341_a;
  wire [32:0] c341_d;
  wire c340_r;
  wire c340_a;
  wire [32:0] c340_d;
  wire c339_r;
  wire c339_a;
  wire [32:0] c339_d;
  wire c338_r;
  wire c338_a;
  wire [32:0] c338_d;
  wire c337_r;
  wire c337_a;
  wire c336_r;
  wire c336_a;
  wire c335_r;
  wire c335_a;
  wire c334_r;
  wire c334_a;
  wire [32:0] c334_d;
  wire c333_r;
  wire c333_a;
  wire [32:0] c333_d;
  wire c332_r;
  wire c332_a;
  wire [31:0] c332_d;
  wire c331_r;
  wire c331_a;
  wire c331_d;
  wire c330_r;
  wire c330_a;
  wire c330_d;
  wire c329_r;
  wire c329_a;
  wire c329_d;
  wire c328_r;
  wire c328_a;
  wire c327_r;
  wire c327_a;
  wire c326_r;
  wire c326_a;
  wire c326_d;
  wire c325_r;
  wire c325_a;
  wire c324_r;
  wire c324_a;
  wire c324_d;
  wire c323_r;
  wire c323_a;
  wire c323_d;
  wire c322_r;
  wire c322_a;
  wire c322_d;
  wire c321_r;
  wire c321_a;
  wire c321_d;
  wire c320_r;
  wire c320_a;
  wire c320_d;
  wire c319_r;
  wire c319_a;
  wire [32:0] c319_d;
  wire c318_r;
  wire c318_a;
  wire [32:0] c318_d;
  wire c317_r;
  wire c317_a;
  wire c316_r;
  wire c316_a;
  wire c315_r;
  wire c315_a;
  wire c314_r;
  wire c314_a;
  wire [32:0] c314_d;
  wire c313_r;
  wire c313_a;
  wire [32:0] c313_d;
  wire c312_r;
  wire c312_a;
  wire [31:0] c312_d;
  wire c311_r;
  wire c311_a;
  wire [33:0] c311_d;
  wire c310_r;
  wire c310_a;
  wire [32:0] c310_d;
  wire c309_r;
  wire c309_a;
  wire [32:0] c309_d;
  wire c308_r;
  wire c308_a;
  wire c308_d;
  wire c307_r;
  wire c307_a;
  wire [33:0] c307_d;
  wire c306_r;
  wire c306_a;
  wire [32:0] c306_d;
  wire c305_r;
  wire c305_a;
  wire [32:0] c305_d;
  wire c304_r;
  wire c304_a;
  wire c304_d;
  wire c303_r;
  wire c303_a;
  wire c303_d;
  wire c302_r;
  wire c302_a;
  wire c302_d;
  wire c301_r;
  wire c301_a;
  wire c301_d;
  wire c300_r;
  wire c300_a;
  wire [32:0] c300_d;
  wire c299_r;
  wire c299_a;
  wire [32:0] c299_d;
  wire c298_r;
  wire c298_a;
  wire c297_r;
  wire c297_a;
  wire c296_r;
  wire c296_a;
  wire c295_r;
  wire c295_a;
  wire [32:0] c295_d;
  wire c294_r;
  wire c294_a;
  wire [32:0] c294_d;
  wire c293_r;
  wire c293_a;
  wire [31:0] c293_d;
  wire c292_r;
  wire c292_a;
  wire [33:0] c292_d;
  wire c291_r;
  wire c291_a;
  wire [32:0] c291_d;
  wire c290_r;
  wire c290_a;
  wire [32:0] c290_d;
  wire c289_r;
  wire c289_a;
  wire c289_d;
  wire c288_r;
  wire c288_a;
  wire [33:0] c288_d;
  wire c287_r;
  wire c287_a;
  wire [32:0] c287_d;
  wire c286_r;
  wire c286_a;
  wire [32:0] c286_d;
  wire c285_r;
  wire c285_a;
  wire [32:0] c285_d;
  wire c284_r;
  wire c284_a;
  wire [32:0] c284_d;
  wire c283_r;
  wire c283_a;
  wire c282_r;
  wire c282_a;
  wire c281_r;
  wire c281_a;
  wire c280_r;
  wire c280_a;
  wire [32:0] c280_d;
  wire c279_r;
  wire c279_a;
  wire [32:0] c279_d;
  wire c278_r;
  wire c278_a;
  wire [31:0] c278_d;
  wire c277_r;
  wire c277_a;
  wire c277_d;
  wire c276_r;
  wire c276_a;
  wire c276_d;
  wire c275_r;
  wire c275_a;
  wire c275_d;
  wire c274_r;
  wire c274_a;
  wire c273_r;
  wire c273_a;
  wire c272_r;
  wire c272_a;
  wire c272_d;
  wire c271_r;
  wire c271_a;
  wire c270_r;
  wire c270_a;
  wire c270_d;
  wire c269_r;
  wire c269_a;
  wire c269_d;
  wire c268_r;
  wire c268_a;
  wire c268_d;
  wire c267_r;
  wire c267_a;
  wire c267_d;
  wire c266_r;
  wire c266_a;
  wire c266_d;
  wire c265_r;
  wire c265_a;
  wire [32:0] c265_d;
  wire c264_r;
  wire c264_a;
  wire [32:0] c264_d;
  wire c263_r;
  wire c263_a;
  wire c262_r;
  wire c262_a;
  wire c261_r;
  wire c261_a;
  wire c260_r;
  wire c260_a;
  wire [32:0] c260_d;
  wire c259_r;
  wire c259_a;
  wire [32:0] c259_d;
  wire c258_r;
  wire c258_a;
  wire [31:0] c258_d;
  wire c257_r;
  wire c257_a;
  wire [33:0] c257_d;
  wire c256_r;
  wire c256_a;
  wire [32:0] c256_d;
  wire c255_r;
  wire c255_a;
  wire [32:0] c255_d;
  wire c254_r;
  wire c254_a;
  wire c254_d;
  wire c253_r;
  wire c253_a;
  wire [33:0] c253_d;
  wire c252_r;
  wire c252_a;
  wire [32:0] c252_d;
  wire c251_r;
  wire c251_a;
  wire [32:0] c251_d;
  wire c250_r;
  wire c250_a;
  wire c250_d;
  wire c249_r;
  wire c249_a;
  wire c249_d;
  wire c248_r;
  wire c248_a;
  wire c248_d;
  wire c247_r;
  wire c247_a;
  wire c247_d;
  wire c246_r;
  wire c246_a;
  wire [32:0] c246_d;
  wire c245_r;
  wire c245_a;
  wire [32:0] c245_d;
  wire c244_r;
  wire c244_a;
  wire c243_r;
  wire c243_a;
  wire c242_r;
  wire c242_a;
  wire c241_r;
  wire c241_a;
  wire [32:0] c241_d;
  wire c240_r;
  wire c240_a;
  wire [32:0] c240_d;
  wire c239_r;
  wire c239_a;
  wire [31:0] c239_d;
  wire c238_r;
  wire c238_a;
  wire [33:0] c238_d;
  wire c237_r;
  wire c237_a;
  wire [32:0] c237_d;
  wire c236_r;
  wire c236_a;
  wire [32:0] c236_d;
  wire c235_r;
  wire c235_a;
  wire c235_d;
  wire c234_r;
  wire c234_a;
  wire [33:0] c234_d;
  wire c233_r;
  wire c233_a;
  wire [32:0] c233_d;
  wire c232_r;
  wire c232_a;
  wire [32:0] c232_d;
  wire c231_r;
  wire c231_a;
  wire [32:0] c231_d;
  wire c230_r;
  wire c230_a;
  wire [32:0] c230_d;
  wire c229_r;
  wire c229_a;
  wire c228_r;
  wire c228_a;
  wire c227_r;
  wire c227_a;
  wire c226_r;
  wire c226_a;
  wire [32:0] c226_d;
  wire c225_r;
  wire c225_a;
  wire [32:0] c225_d;
  wire c224_r;
  wire c224_a;
  wire [31:0] c224_d;
  wire c223_r;
  wire c223_a;
  wire c223_d;
  wire c222_r;
  wire c222_a;
  wire c222_d;
  wire c221_r;
  wire c221_a;
  wire c221_d;
  wire c220_r;
  wire c220_a;
  wire c219_r;
  wire c219_a;
  wire c218_r;
  wire c218_a;
  wire c218_d;
  wire c217_r;
  wire c217_a;
  wire c216_r;
  wire c216_a;
  wire c216_d;
  wire c215_r;
  wire c215_a;
  wire c215_d;
  wire c214_r;
  wire c214_a;
  wire c214_d;
  wire c213_r;
  wire c213_a;
  wire c213_d;
  wire c212_r;
  wire c212_a;
  wire c212_d;
  wire c211_r;
  wire c211_a;
  wire [32:0] c211_d;
  wire c210_r;
  wire c210_a;
  wire [32:0] c210_d;
  wire c209_r;
  wire c209_a;
  wire c208_r;
  wire c208_a;
  wire c207_r;
  wire c207_a;
  wire c206_r;
  wire c206_a;
  wire [32:0] c206_d;
  wire c205_r;
  wire c205_a;
  wire [32:0] c205_d;
  wire c204_r;
  wire c204_a;
  wire [31:0] c204_d;
  wire c203_r;
  wire c203_a;
  wire [33:0] c203_d;
  wire c202_r;
  wire c202_a;
  wire [32:0] c202_d;
  wire c201_r;
  wire c201_a;
  wire [32:0] c201_d;
  wire c200_r;
  wire c200_a;
  wire c200_d;
  wire c199_r;
  wire c199_a;
  wire [33:0] c199_d;
  wire c198_r;
  wire c198_a;
  wire [32:0] c198_d;
  wire c197_r;
  wire c197_a;
  wire [32:0] c197_d;
  wire c196_r;
  wire c196_a;
  wire c196_d;
  wire c195_r;
  wire c195_a;
  wire c195_d;
  wire c194_r;
  wire c194_a;
  wire c194_d;
  wire c193_r;
  wire c193_a;
  wire c193_d;
  wire c192_r;
  wire c192_a;
  wire [32:0] c192_d;
  wire c191_r;
  wire c191_a;
  wire [32:0] c191_d;
  wire c190_r;
  wire c190_a;
  wire c189_r;
  wire c189_a;
  wire c188_r;
  wire c188_a;
  wire c187_r;
  wire c187_a;
  wire [32:0] c187_d;
  wire c186_r;
  wire c186_a;
  wire [32:0] c186_d;
  wire c185_r;
  wire c185_a;
  wire [31:0] c185_d;
  wire c184_r;
  wire c184_a;
  wire [33:0] c184_d;
  wire c183_r;
  wire c183_a;
  wire [32:0] c183_d;
  wire c182_r;
  wire c182_a;
  wire [32:0] c182_d;
  wire c181_r;
  wire c181_a;
  wire c181_d;
  wire c180_r;
  wire c180_a;
  wire [33:0] c180_d;
  wire c179_r;
  wire c179_a;
  wire [32:0] c179_d;
  wire c178_r;
  wire c178_a;
  wire [32:0] c178_d;
  wire c177_r;
  wire c177_a;
  wire [32:0] c177_d;
  wire c176_r;
  wire c176_a;
  wire [32:0] c176_d;
  wire c175_r;
  wire c175_a;
  wire c174_r;
  wire c174_a;
  wire c173_r;
  wire c173_a;
  wire c172_r;
  wire c172_a;
  wire [32:0] c172_d;
  wire c171_r;
  wire c171_a;
  wire [32:0] c171_d;
  wire c170_r;
  wire c170_a;
  wire [31:0] c170_d;
  wire c169_r;
  wire c169_a;
  wire c169_d;
  wire c168_r;
  wire c168_a;
  wire c168_d;
  wire c167_r;
  wire c167_a;
  wire c167_d;
  wire c166_r;
  wire c166_a;
  wire c165_r;
  wire c165_a;
  wire c164_r;
  wire c164_a;
  wire c164_d;
  wire c163_r;
  wire c163_a;
  wire c162_r;
  wire c162_a;
  wire c162_d;
  wire c161_r;
  wire c161_a;
  wire c161_d;
  wire c160_r;
  wire c160_a;
  wire c160_d;
  wire c159_r;
  wire c159_a;
  wire c159_d;
  wire c158_r;
  wire c158_a;
  wire c158_d;
  wire c157_r;
  wire c157_a;
  wire [32:0] c157_d;
  wire c156_r;
  wire c156_a;
  wire [32:0] c156_d;
  wire c155_r;
  wire c155_a;
  wire c154_r;
  wire c154_a;
  wire c153_r;
  wire c153_a;
  wire c152_r;
  wire c152_a;
  wire [32:0] c152_d;
  wire c151_r;
  wire c151_a;
  wire [32:0] c151_d;
  wire c150_r;
  wire c150_a;
  wire [31:0] c150_d;
  wire c149_r;
  wire c149_a;
  wire [33:0] c149_d;
  wire c148_r;
  wire c148_a;
  wire [32:0] c148_d;
  wire c147_r;
  wire c147_a;
  wire [32:0] c147_d;
  wire c146_r;
  wire c146_a;
  wire c146_d;
  wire c145_r;
  wire c145_a;
  wire [33:0] c145_d;
  wire c144_r;
  wire c144_a;
  wire [32:0] c144_d;
  wire c143_r;
  wire c143_a;
  wire [32:0] c143_d;
  wire c142_r;
  wire c142_a;
  wire c142_d;
  wire c141_r;
  wire c141_a;
  wire c141_d;
  wire c140_r;
  wire c140_a;
  wire c140_d;
  wire c139_r;
  wire c139_a;
  wire c139_d;
  wire c138_r;
  wire c138_a;
  wire [32:0] c138_d;
  wire c137_r;
  wire c137_a;
  wire [32:0] c137_d;
  wire c136_r;
  wire c136_a;
  wire c135_r;
  wire c135_a;
  wire c134_r;
  wire c134_a;
  wire c133_r;
  wire c133_a;
  wire [32:0] c133_d;
  wire c132_r;
  wire c132_a;
  wire [32:0] c132_d;
  wire c131_r;
  wire c131_a;
  wire [31:0] c131_d;
  wire c130_r;
  wire c130_a;
  wire [33:0] c130_d;
  wire c129_r;
  wire c129_a;
  wire [32:0] c129_d;
  wire c128_r;
  wire c128_a;
  wire [32:0] c128_d;
  wire c127_r;
  wire c127_a;
  wire c127_d;
  wire c126_r;
  wire c126_a;
  wire [33:0] c126_d;
  wire c125_r;
  wire c125_a;
  wire [32:0] c125_d;
  wire c124_r;
  wire c124_a;
  wire [32:0] c124_d;
  wire c123_r;
  wire c123_a;
  wire [32:0] c123_d;
  wire c122_r;
  wire c122_a;
  wire [32:0] c122_d;
  wire c121_r;
  wire c121_a;
  wire c120_r;
  wire c120_a;
  wire c119_r;
  wire c119_a;
  wire c118_r;
  wire c118_a;
  wire [32:0] c118_d;
  wire c117_r;
  wire c117_a;
  wire [32:0] c117_d;
  wire c116_r;
  wire c116_a;
  wire [31:0] c116_d;
  wire c115_r;
  wire c115_a;
  wire c115_d;
  wire c114_r;
  wire c114_a;
  wire c114_d;
  wire c113_r;
  wire c113_a;
  wire c113_d;
  wire c112_r;
  wire c112_a;
  wire c111_r;
  wire c111_a;
  wire c110_r;
  wire c110_a;
  wire c110_d;
  wire c109_r;
  wire c109_a;
  wire c108_r;
  wire c108_a;
  wire c108_d;
  wire c107_r;
  wire c107_a;
  wire c107_d;
  wire c106_r;
  wire c106_a;
  wire c106_d;
  wire c105_r;
  wire c105_a;
  wire c105_d;
  wire c104_r;
  wire c104_a;
  wire c104_d;
  wire c103_r;
  wire c103_a;
  wire [32:0] c103_d;
  wire c102_r;
  wire c102_a;
  wire [32:0] c102_d;
  wire c101_r;
  wire c101_a;
  wire c100_r;
  wire c100_a;
  wire c99_r;
  wire c99_a;
  wire c98_r;
  wire c98_a;
  wire [32:0] c98_d;
  wire c97_r;
  wire c97_a;
  wire [32:0] c97_d;
  wire c96_r;
  wire c96_a;
  wire [31:0] c96_d;
  wire c95_r;
  wire c95_a;
  wire [33:0] c95_d;
  wire c94_r;
  wire c94_a;
  wire [32:0] c94_d;
  wire c93_r;
  wire c93_a;
  wire [32:0] c93_d;
  wire c92_r;
  wire c92_a;
  wire c92_d;
  wire c91_r;
  wire c91_a;
  wire [33:0] c91_d;
  wire c90_r;
  wire c90_a;
  wire [32:0] c90_d;
  wire c89_r;
  wire c89_a;
  wire [32:0] c89_d;
  wire c88_r;
  wire c88_a;
  wire c88_d;
  wire c87_r;
  wire c87_a;
  wire c87_d;
  wire c86_r;
  wire c86_a;
  wire c86_d;
  wire c85_r;
  wire c85_a;
  wire c85_d;
  wire c84_r;
  wire c84_a;
  wire [32:0] c84_d;
  wire c83_r;
  wire c83_a;
  wire [32:0] c83_d;
  wire c82_r;
  wire c82_a;
  wire c81_r;
  wire c81_a;
  wire c80_r;
  wire c80_a;
  wire c79_r;
  wire c79_a;
  wire [32:0] c79_d;
  wire c78_r;
  wire c78_a;
  wire [32:0] c78_d;
  wire c77_r;
  wire c77_a;
  wire [31:0] c77_d;
  wire c76_r;
  wire c76_a;
  wire [33:0] c76_d;
  wire c75_r;
  wire c75_a;
  wire [32:0] c75_d;
  wire c74_r;
  wire c74_a;
  wire [32:0] c74_d;
  wire c73_r;
  wire c73_a;
  wire c73_d;
  wire c72_r;
  wire c72_a;
  wire [33:0] c72_d;
  wire c71_r;
  wire c71_a;
  wire [32:0] c71_d;
  wire c70_r;
  wire c70_a;
  wire [32:0] c70_d;
  wire c69_r;
  wire c69_a;
  wire [32:0] c69_d;
  wire c68_r;
  wire c68_a;
  wire [32:0] c68_d;
  wire c67_r;
  wire c67_a;
  wire c66_r;
  wire c66_a;
  wire c65_r;
  wire c65_a;
  wire c64_r;
  wire c64_a;
  wire [32:0] c64_d;
  wire c63_r;
  wire c63_a;
  wire [32:0] c63_d;
  wire c62_r;
  wire c62_a;
  wire [31:0] c62_d;
  wire c61_r;
  wire c61_a;
  wire c61_d;
  wire c60_r;
  wire c60_a;
  wire c60_d;
  wire c59_r;
  wire c59_a;
  wire c59_d;
  wire c58_r;
  wire c58_a;
  wire c57_r;
  wire c57_a;
  wire c56_r;
  wire c56_a;
  wire c56_d;
  wire c55_r;
  wire c55_a;
  wire c54_r;
  wire c54_a;
  wire c54_d;
  wire c53_r;
  wire c53_a;
  wire c53_d;
  wire c52_r;
  wire c52_a;
  wire c52_d;
  wire c51_r;
  wire c51_a;
  wire c51_d;
  wire c50_r;
  wire c50_a;
  wire c50_d;
  wire c49_r;
  wire c49_a;
  wire [32:0] c49_d;
  wire c48_r;
  wire c48_a;
  wire [32:0] c48_d;
  wire c47_r;
  wire c47_a;
  wire c46_r;
  wire c46_a;
  wire c45_r;
  wire c45_a;
  wire c44_r;
  wire c44_a;
  wire [32:0] c44_d;
  wire c43_r;
  wire c43_a;
  wire [32:0] c43_d;
  wire c42_r;
  wire c42_a;
  wire [31:0] c42_d;
  wire c41_r;
  wire c41_a;
  wire [33:0] c41_d;
  wire c40_r;
  wire c40_a;
  wire [32:0] c40_d;
  wire c39_r;
  wire c39_a;
  wire [32:0] c39_d;
  wire c38_r;
  wire c38_a;
  wire c38_d;
  wire c37_r;
  wire c37_a;
  wire [33:0] c37_d;
  wire c36_r;
  wire c36_a;
  wire [32:0] c36_d;
  wire c35_r;
  wire c35_a;
  wire [32:0] c35_d;
  wire c34_r;
  wire c34_a;
  wire c34_d;
  wire c33_r;
  wire c33_a;
  wire c33_d;
  wire c32_r;
  wire c32_a;
  wire c32_d;
  wire c31_r;
  wire c31_a;
  wire c31_d;
  wire c30_r;
  wire c30_a;
  wire [32:0] c30_d;
  wire c29_r;
  wire c29_a;
  wire [32:0] c29_d;
  wire c28_r;
  wire c28_a;
  wire c27_r;
  wire c27_a;
  wire c26_r;
  wire c26_a;
  wire c25_r;
  wire c25_a;
  wire [32:0] c25_d;
  wire c24_r;
  wire c24_a;
  wire [32:0] c24_d;
  wire c23_r;
  wire c23_a;
  wire [31:0] c23_d;
  wire c22_r;
  wire c22_a;
  wire [33:0] c22_d;
  wire c21_r;
  wire c21_a;
  wire [32:0] c21_d;
  wire c20_r;
  wire c20_a;
  wire [32:0] c20_d;
  wire c19_r;
  wire c19_a;
  wire c19_d;
  wire c18_r;
  wire c18_a;
  wire [33:0] c18_d;
  wire c17_r;
  wire c17_a;
  wire [32:0] c17_d;
  wire c16_r;
  wire c16_a;
  wire [32:0] c16_d;
  wire c15_r;
  wire c15_a;
  wire [32:0] c15_d;
  wire c14_r;
  wire c14_a;
  wire [32:0] c14_d;
  wire c13_r;
  wire c13_a;
  wire c12_r;
  wire c12_a;
  wire c11_r;
  wire c11_a;
  wire c10_r;
  wire c10_a;
  wire [32:0] c10_d;
  wire c9_r;
  wire c9_a;
  wire [32:0] c9_d;
  wire c8_r;
  wire c8_a;
  wire [31:0] c8_d;
  wire c7_r;
  wire c7_a;
  wire c7_d;
  wire c6_r;
  wire c6_a;
  wire c5_r;
  wire c5_a;
  wire [31:0] c5_d;
  BrzVariable_16_2_s0_ I0 (c891_r, c891_a, c891_d, c883_r, c883_a, c883_d, c877_r, c877_a, c877_d);
  BrzVariable_16_1_s0_ I1 (c889_r, c889_a, c889_d, c871_r, c871_a, c871_d);
  BrzVariable_33_32_s0_ I2 (c886_r, c886_a, c886_d, c830_r, c830_a, c830_d, c826_r, c826_a, c826_d, c776_r, c776_a, c776_d, c772_r, c772_a, c772_d, c722_r, c722_a, c722_d, c718_r, c718_a, c718_d, c668_r, c668_a, c668_d, c664_r, c664_a, c664_d, c614_r, c614_a, c614_d, c610_r, c610_a, c610_d, c560_r, c560_a, c560_d, c556_r, c556_a, c556_d, c506_r, c506_a, c506_d, c502_r, c502_a, c502_d, c452_r, c452_a, c452_d, c448_r, c448_a,
		c448_d, c398_r, c398_a, c398_d, c394_r, c394_a, c394_d, c344_r, c344_a, c344_d, c340_r, c340_a, c340_d, c290_r, c290_a, c290_d, c286_r, c286_a, c286_d, c236_r, c236_a, c236_d, c232_r, c232_a, c232_d, c182_r, c182_a, c182_d, c178_r, c178_a, c178_d, c128_r, c128_a, c128_d, c124_r, c124_a, c124_d, c74_r, c74_a, c74_d, c70_r, c70_a, c70_d, c20_r, c20_a, c20_d, c16_r, c16_a, c16_d);
  BrzVariable_33_32_s0_ I3 (c881_r, c881_a, c881_d, c849_r, c849_a, c849_d, c845_r, c845_a, c845_d, c795_r, c795_a, c795_d, c791_r, c791_a, c791_d, c741_r, c741_a, c741_d, c737_r, c737_a, c737_d, c687_r, c687_a, c687_d, c683_r, c683_a, c683_d, c633_r, c633_a, c633_d, c629_r, c629_a, c629_d, c579_r, c579_a, c579_d, c575_r, c575_a, c575_d, c525_r, c525_a, c525_d, c521_r, c521_a, c521_d, c471_r, c471_a, c471_d, c467_r, c467_a,
		c467_d, c417_r, c417_a, c417_d, c413_r, c413_a, c413_d, c363_r, c363_a, c363_d, c359_r, c359_a, c359_d, c309_r, c309_a, c309_d, c305_r, c305_a, c305_d, c255_r, c255_a, c255_d, c251_r, c251_a, c251_d, c201_r, c201_a, c201_d, c197_r, c197_a, c197_d, c147_r, c147_a, c147_d, c143_r, c143_a, c143_d, c93_r, c93_a, c93_d, c89_r, c89_a, c89_d, c39_r, c39_a, c39_d, c35_r, c35_a, c35_d);
  BrzVariable_33_161_s1305_1_2e_2e1_3b0_2e_2_m4m I4 (c895_r, c895_a, c895_d, c862_r, c862_a, c862_d, c860_r, c860_a, c860_d, c842_r, c842_a, c842_d, c841_r, c841_a, c841_d, c850_r, c850_a, c850_d, c846_r, c846_a, c846_d, c831_r, c831_a, c831_d, c827_r, c827_a, c827_d, c818_r, c818_a, c818_d, c817_r, c817_a, c817_d, c808_r, c808_a, c808_d, c806_r, c806_a, c806_d, c788_r, c788_a, c788_d, c787_r, c787_a, c787_d, c796_r, c796_a, c796_d, c792_r, c792_a,
		c792_d, c777_r, c777_a, c777_d, c773_r, c773_a, c773_d, c764_r, c764_a, c764_d, c763_r, c763_a, c763_d, c754_r, c754_a, c754_d, c752_r, c752_a, c752_d, c734_r, c734_a, c734_d, c733_r, c733_a, c733_d, c742_r, c742_a, c742_d, c738_r, c738_a, c738_d, c723_r, c723_a, c723_d, c719_r, c719_a, c719_d, c710_r, c710_a, c710_d, c709_r, c709_a, c709_d, c700_r, c700_a, c700_d, c698_r, c698_a, c698_d, c680_r, c680_a,
		c680_d, c679_r, c679_a, c679_d, c688_r, c688_a, c688_d, c684_r, c684_a, c684_d, c669_r, c669_a, c669_d, c665_r, c665_a, c665_d, c656_r, c656_a, c656_d, c655_r, c655_a, c655_d, c646_r, c646_a, c646_d, c644_r, c644_a, c644_d, c626_r, c626_a, c626_d, c625_r, c625_a, c625_d, c634_r, c634_a, c634_d, c630_r, c630_a, c630_d, c615_r, c615_a, c615_d, c611_r, c611_a, c611_d, c602_r, c602_a, c602_d, c601_r, c601_a,
		c601_d, c592_r, c592_a, c592_d, c590_r, c590_a, c590_d, c572_r, c572_a, c572_d, c571_r, c571_a, c571_d, c580_r, c580_a, c580_d, c576_r, c576_a, c576_d, c561_r, c561_a, c561_d, c557_r, c557_a, c557_d, c548_r, c548_a, c548_d, c547_r, c547_a, c547_d, c538_r, c538_a, c538_d, c536_r, c536_a, c536_d, c518_r, c518_a, c518_d, c517_r, c517_a, c517_d, c526_r, c526_a, c526_d, c522_r, c522_a, c522_d, c507_r, c507_a,
		c507_d, c503_r, c503_a, c503_d, c494_r, c494_a, c494_d, c493_r, c493_a, c493_d, c484_r, c484_a, c484_d, c482_r, c482_a, c482_d, c464_r, c464_a, c464_d, c463_r, c463_a, c463_d, c472_r, c472_a, c472_d, c468_r, c468_a, c468_d, c453_r, c453_a, c453_d, c449_r, c449_a, c449_d, c440_r, c440_a, c440_d, c439_r, c439_a, c439_d, c430_r, c430_a, c430_d, c428_r, c428_a, c428_d, c410_r, c410_a, c410_d, c409_r, c409_a,
		c409_d, c418_r, c418_a, c418_d, c414_r, c414_a, c414_d, c399_r, c399_a, c399_d, c395_r, c395_a, c395_d, c386_r, c386_a, c386_d, c385_r, c385_a, c385_d, c376_r, c376_a, c376_d, c374_r, c374_a, c374_d, c356_r, c356_a, c356_d, c355_r, c355_a, c355_d, c364_r, c364_a, c364_d, c360_r, c360_a, c360_d, c345_r, c345_a, c345_d, c341_r, c341_a, c341_d, c332_r, c332_a, c332_d, c331_r, c331_a, c331_d, c322_r, c322_a,
		c322_d, c320_r, c320_a, c320_d, c302_r, c302_a, c302_d, c301_r, c301_a, c301_d, c310_r, c310_a, c310_d, c306_r, c306_a, c306_d, c291_r, c291_a, c291_d, c287_r, c287_a, c287_d, c278_r, c278_a, c278_d, c277_r, c277_a, c277_d, c268_r, c268_a, c268_d, c266_r, c266_a, c266_d, c248_r, c248_a, c248_d, c247_r, c247_a, c247_d, c256_r, c256_a, c256_d, c252_r, c252_a, c252_d, c237_r, c237_a, c237_d, c233_r, c233_a,
		c233_d, c224_r, c224_a, c224_d, c223_r, c223_a, c223_d, c214_r, c214_a, c214_d, c212_r, c212_a, c212_d, c194_r, c194_a, c194_d, c193_r, c193_a, c193_d, c202_r, c202_a, c202_d, c198_r, c198_a, c198_d, c183_r, c183_a, c183_d, c179_r, c179_a, c179_d, c170_r, c170_a, c170_d, c169_r, c169_a, c169_d, c160_r, c160_a, c160_d, c158_r, c158_a, c158_d, c140_r, c140_a, c140_d, c139_r, c139_a, c139_d, c148_r, c148_a,
		c148_d, c144_r, c144_a, c144_d, c129_r, c129_a, c129_d, c125_r, c125_a, c125_d, c116_r, c116_a, c116_d, c115_r, c115_a, c115_d, c106_r, c106_a, c106_d, c104_r, c104_a, c104_d, c86_r, c86_a, c86_d, c85_r, c85_a, c85_d, c94_r, c94_a, c94_d, c90_r, c90_a, c90_d, c75_r, c75_a, c75_d, c71_r, c71_a, c71_d, c62_r, c62_a, c62_d, c61_r, c61_a, c61_d, c52_r, c52_a, c52_d, c50_r, c50_a,
		c50_d, c32_r, c32_a, c32_d, c31_r, c31_a, c31_d, c40_r, c40_a, c40_d, c36_r, c36_a, c36_d, c21_r, c21_a, c21_d, c17_r, c17_a, c17_d, c8_r, c8_a, c8_d, c7_r, c7_a, c7_d, c5_r, c5_a, c5_d);
  BrzCallMux_33_49 I5 (c10_r, c10_a, c10_d, c25_r, c25_a, c25_d, c44_r, c44_a, c44_d, c64_r, c64_a, c64_d, c79_r, c79_a, c79_d, c98_r, c98_a, c98_d, c118_r, c118_a, c118_d, c133_r, c133_a, c133_d, c152_r, c152_a, c152_d, c172_r, c172_a, c172_d, c187_r, c187_a, c187_d, c206_r, c206_a, c206_d, c226_r, c226_a, c226_d, c241_r, c241_a, c241_d, c260_r, c260_a, c260_d, c280_r, c280_a, c280_d, c295_r, c295_a,
		c295_d, c314_r, c314_a, c314_d, c334_r, c334_a, c334_d, c349_r, c349_a, c349_d, c368_r, c368_a, c368_d, c388_r, c388_a, c388_d, c403_r, c403_a, c403_d, c422_r, c422_a, c422_d, c442_r, c442_a, c442_d, c457_r, c457_a, c457_d, c476_r, c476_a, c476_d, c496_r, c496_a, c496_d, c511_r, c511_a, c511_d, c530_r, c530_a, c530_d, c550_r, c550_a, c550_d, c565_r, c565_a, c565_d, c584_r, c584_a, c584_d, c604_r, c604_a,
		c604_d, c619_r, c619_a, c619_d, c638_r, c638_a, c638_d, c658_r, c658_a, c658_d, c673_r, c673_a, c673_d, c692_r, c692_a, c692_d, c712_r, c712_a, c712_d, c727_r, c727_a, c727_d, c746_r, c746_a, c746_d, c766_r, c766_a, c766_d, c781_r, c781_a, c781_d, c800_r, c800_a, c800_d, c820_r, c820_a, c820_d, c835_r, c835_a, c835_d, c854_r, c854_a, c854_d, c875_r, c875_a, c875_d, c895_r, c895_a, c895_d);
  BrzLoop I6 (activate_0r, activate_0a, c894_r, c894_a);
  BrzSequence_35_s34_SSSSSSSSSSSSSSSSSSSSSSS_m3m I7 (c894_r, c894_a, c893_r, c893_a, c888_r, c888_a, c867_r, c867_a, c868_r, c868_a, c813_r, c813_a, c814_r, c814_a, c759_r, c759_a, c760_r, c760_a, c705_r, c705_a, c706_r, c706_a, c651_r, c651_a, c652_r, c652_a, c597_r, c597_a, c598_r, c598_a, c543_r, c543_a, c544_r, c544_a, c489_r, c489_a, c490_r, c490_a, c435_r, c435_a, c436_r, c436_a, c381_r, c381_a, c382_r, c382_a, c327_r, c327_a, c328_r, c328_a,
		c273_r, c273_a, c274_r, c274_a, c219_r, c219_a, c220_r, c220_a, c165_r, c165_a, c166_r, c166_a, c111_r, c111_a, c112_r, c112_a, c57_r, c57_a, c58_r, c58_a, c6_r, c6_a);
  BrzConcur_2 I8 (c893_r, c893_a, c892_r, c892_a, c890_r, c890_a);
  BrzFetch_16_s5_false I9 (c892_r, c892_a, x_0r, x_0a, x_0d, c891_r, c891_a, c891_d);
  BrzFetch_16_s5_false I10 (c890_r, c890_a, y_0r, y_0a, y_0d, c889_r, c889_a, c889_d);
  BrzConcur_3 I11 (c888_r, c888_a, c887_r, c887_a, c882_r, c882_a, c876_r, c876_a);
  BrzFetch_33_s5_false I12 (c887_r, c887_a, c885_r, c885_a, c885_d, c886_r, c886_a, c886_d);
  BrzCombine_33_17_16 I13 (c885_r, c885_a, c885_d, c884_r, c884_a, c884_d, c883_r, c883_a, c883_d);
  BrzConstant_17_0 I14 (c884_r, c884_a, c884_d);
  BrzFetch_33_s5_false I15 (c882_r, c882_a, c880_r, c880_a, c880_d, c881_r, c881_a, c881_d);
  BrzCombine_33_17_16 I16 (c880_r, c880_a, c880_d, c879_r, c879_a, c879_d, c878_r, c878_a, c878_d);
  BrzConstant_17_0 I17 (c879_r, c879_a, c879_d);
  BrzUnaryFunc_16_16_s6_Negate_s4_true I18 (c878_r, c878_a, c878_d, c877_r, c877_a, c877_d);
  BrzFetch_33_s5_false I19 (c876_r, c876_a, c874_r, c874_a, c874_d, c875_r, c875_a, c875_d);
  BrzAdapt_33_17_s5_false_s5_false I20 (c874_r, c874_a, c874_d, c873_r, c873_a, c873_d);
  BrzCombine_17_1_16 I21 (c873_r, c873_a, c873_d, c872_r, c872_a, c872_d, c871_r, c871_a, c871_d);
  BrzConstant_1_0 I22 (c872_r, c872_a, c872_d);
  BrzCase_1_2_s5_0_3b1 I23 (c866_r, c866_a, c866_d, c821_r, c821_a, c865_r, c865_a);
  BrzFetch_1_s5_false I24 (c867_r, c867_a, c864_r, c864_a, c864_d, c869_r, c869_a, c869_d);
  BrzFetch_1_s5_false I25 (c868_r, c868_a, c870_r, c870_a, c870_d, c866_r, c866_a, c866_d);
  BrzVariable_1_1_s0_ I26 (c869_r, c869_a, c869_d, c870_r, c870_a, c870_d);
  BrzBar_2 I27 (c864_r, c864_a, c864_d, c865_r, c865_a, c844_r, c844_a, c844_d, c863_r, c863_a, c863_d, c836_r, c836_a, c855_r, c855_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I28 (c863_r, c863_a, c863_d, c862_r, c862_a, c862_d, c861_r, c861_a, c861_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I29 (c861_r, c861_a, c861_d, c860_r, c860_a, c860_d);
  BrzSequence_2_s1_S I30 (c855_r, c855_a, c856_r, c856_a, c857_r, c857_a);
  BrzFetch_33_s5_false I31 (c856_r, c856_a, c853_r, c853_a, c853_d, c858_r, c858_a, c858_d);
  BrzFetch_33_s5_false I32 (c857_r, c857_a, c859_r, c859_a, c859_d, c854_r, c854_a, c854_d);
  BrzVariable_33_1_s0_ I33 (c858_r, c858_a, c858_d, c859_r, c859_a, c859_d);
  BrzCombine_33_32_1 I34 (c853_r, c853_a, c853_d, c852_r, c852_a, c852_d, c848_r, c848_a, c848_d);
  BrzSlice_32_34_1 I35 (c852_r, c852_a, c852_d, c851_r, c851_a, c851_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I36 (c851_r, c851_a, c851_d, c850_r, c850_a, c850_d, c849_r, c849_a, c849_d);
  BrzSlice_1_34_32 I37 (c848_r, c848_a, c848_d, c847_r, c847_a, c847_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I38 (c847_r, c847_a, c847_d, c846_r, c846_a, c846_d, c845_r, c845_a, c845_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I39 (c844_r, c844_a, c844_d, c843_r, c843_a, c843_d, c841_r, c841_a, c841_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I40 (c843_r, c843_a, c843_d, c842_r, c842_a, c842_d);
  BrzSequence_2_s1_S I41 (c836_r, c836_a, c837_r, c837_a, c838_r, c838_a);
  BrzFetch_33_s5_false I42 (c837_r, c837_a, c834_r, c834_a, c834_d, c839_r, c839_a, c839_d);
  BrzFetch_33_s5_false I43 (c838_r, c838_a, c840_r, c840_a, c840_d, c835_r, c835_a, c835_d);
  BrzVariable_33_1_s0_ I44 (c839_r, c839_a, c839_d, c840_r, c840_a, c840_d);
  BrzCombine_33_32_1 I45 (c834_r, c834_a, c834_d, c833_r, c833_a, c833_d, c829_r, c829_a, c829_d);
  BrzSlice_32_34_1 I46 (c833_r, c833_a, c833_d, c832_r, c832_a, c832_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I47 (c832_r, c832_a, c832_d, c831_r, c831_a, c831_d, c830_r, c830_a, c830_d);
  BrzSlice_1_34_32 I48 (c829_r, c829_a, c829_d, c828_r, c828_a, c828_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I49 (c828_r, c828_a, c828_d, c827_r, c827_a, c827_d, c826_r, c826_a, c826_d);
  BrzSequence_2_s1_S I50 (c821_r, c821_a, c822_r, c822_a, c823_r, c823_a);
  BrzFetch_33_s5_false I51 (c822_r, c822_a, c819_r, c819_a, c819_d, c824_r, c824_a, c824_d);
  BrzFetch_33_s5_false I52 (c823_r, c823_a, c825_r, c825_a, c825_d, c820_r, c820_a, c820_d);
  BrzVariable_33_1_s0_ I53 (c824_r, c824_a, c824_d, c825_r, c825_a, c825_d);
  BrzCombine_33_32_1 I54 (c819_r, c819_a, c819_d, c818_r, c818_a, c818_d, c817_r, c817_a, c817_d);
  BrzCase_1_2_s5_0_3b1 I55 (c812_r, c812_a, c812_d, c767_r, c767_a, c811_r, c811_a);
  BrzFetch_1_s5_false I56 (c813_r, c813_a, c810_r, c810_a, c810_d, c815_r, c815_a, c815_d);
  BrzFetch_1_s5_false I57 (c814_r, c814_a, c816_r, c816_a, c816_d, c812_r, c812_a, c812_d);
  BrzVariable_1_1_s0_ I58 (c815_r, c815_a, c815_d, c816_r, c816_a, c816_d);
  BrzBar_2 I59 (c810_r, c810_a, c810_d, c811_r, c811_a, c790_r, c790_a, c790_d, c809_r, c809_a, c809_d, c782_r, c782_a, c801_r, c801_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I60 (c809_r, c809_a, c809_d, c808_r, c808_a, c808_d, c807_r, c807_a, c807_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I61 (c807_r, c807_a, c807_d, c806_r, c806_a, c806_d);
  BrzSequence_2_s1_S I62 (c801_r, c801_a, c802_r, c802_a, c803_r, c803_a);
  BrzFetch_33_s5_false I63 (c802_r, c802_a, c799_r, c799_a, c799_d, c804_r, c804_a, c804_d);
  BrzFetch_33_s5_false I64 (c803_r, c803_a, c805_r, c805_a, c805_d, c800_r, c800_a, c800_d);
  BrzVariable_33_1_s0_ I65 (c804_r, c804_a, c804_d, c805_r, c805_a, c805_d);
  BrzCombine_33_32_1 I66 (c799_r, c799_a, c799_d, c798_r, c798_a, c798_d, c794_r, c794_a, c794_d);
  BrzSlice_32_34_1 I67 (c798_r, c798_a, c798_d, c797_r, c797_a, c797_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I68 (c797_r, c797_a, c797_d, c796_r, c796_a, c796_d, c795_r, c795_a, c795_d);
  BrzSlice_1_34_32 I69 (c794_r, c794_a, c794_d, c793_r, c793_a, c793_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I70 (c793_r, c793_a, c793_d, c792_r, c792_a, c792_d, c791_r, c791_a, c791_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I71 (c790_r, c790_a, c790_d, c789_r, c789_a, c789_d, c787_r, c787_a, c787_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I72 (c789_r, c789_a, c789_d, c788_r, c788_a, c788_d);
  BrzSequence_2_s1_S I73 (c782_r, c782_a, c783_r, c783_a, c784_r, c784_a);
  BrzFetch_33_s5_false I74 (c783_r, c783_a, c780_r, c780_a, c780_d, c785_r, c785_a, c785_d);
  BrzFetch_33_s5_false I75 (c784_r, c784_a, c786_r, c786_a, c786_d, c781_r, c781_a, c781_d);
  BrzVariable_33_1_s0_ I76 (c785_r, c785_a, c785_d, c786_r, c786_a, c786_d);
  BrzCombine_33_32_1 I77 (c780_r, c780_a, c780_d, c779_r, c779_a, c779_d, c775_r, c775_a, c775_d);
  BrzSlice_32_34_1 I78 (c779_r, c779_a, c779_d, c778_r, c778_a, c778_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I79 (c778_r, c778_a, c778_d, c777_r, c777_a, c777_d, c776_r, c776_a, c776_d);
  BrzSlice_1_34_32 I80 (c775_r, c775_a, c775_d, c774_r, c774_a, c774_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I81 (c774_r, c774_a, c774_d, c773_r, c773_a, c773_d, c772_r, c772_a, c772_d);
  BrzSequence_2_s1_S I82 (c767_r, c767_a, c768_r, c768_a, c769_r, c769_a);
  BrzFetch_33_s5_false I83 (c768_r, c768_a, c765_r, c765_a, c765_d, c770_r, c770_a, c770_d);
  BrzFetch_33_s5_false I84 (c769_r, c769_a, c771_r, c771_a, c771_d, c766_r, c766_a, c766_d);
  BrzVariable_33_1_s0_ I85 (c770_r, c770_a, c770_d, c771_r, c771_a, c771_d);
  BrzCombine_33_32_1 I86 (c765_r, c765_a, c765_d, c764_r, c764_a, c764_d, c763_r, c763_a, c763_d);
  BrzCase_1_2_s5_0_3b1 I87 (c758_r, c758_a, c758_d, c713_r, c713_a, c757_r, c757_a);
  BrzFetch_1_s5_false I88 (c759_r, c759_a, c756_r, c756_a, c756_d, c761_r, c761_a, c761_d);
  BrzFetch_1_s5_false I89 (c760_r, c760_a, c762_r, c762_a, c762_d, c758_r, c758_a, c758_d);
  BrzVariable_1_1_s0_ I90 (c761_r, c761_a, c761_d, c762_r, c762_a, c762_d);
  BrzBar_2 I91 (c756_r, c756_a, c756_d, c757_r, c757_a, c736_r, c736_a, c736_d, c755_r, c755_a, c755_d, c728_r, c728_a, c747_r, c747_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I92 (c755_r, c755_a, c755_d, c754_r, c754_a, c754_d, c753_r, c753_a, c753_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I93 (c753_r, c753_a, c753_d, c752_r, c752_a, c752_d);
  BrzSequence_2_s1_S I94 (c747_r, c747_a, c748_r, c748_a, c749_r, c749_a);
  BrzFetch_33_s5_false I95 (c748_r, c748_a, c745_r, c745_a, c745_d, c750_r, c750_a, c750_d);
  BrzFetch_33_s5_false I96 (c749_r, c749_a, c751_r, c751_a, c751_d, c746_r, c746_a, c746_d);
  BrzVariable_33_1_s0_ I97 (c750_r, c750_a, c750_d, c751_r, c751_a, c751_d);
  BrzCombine_33_32_1 I98 (c745_r, c745_a, c745_d, c744_r, c744_a, c744_d, c740_r, c740_a, c740_d);
  BrzSlice_32_34_1 I99 (c744_r, c744_a, c744_d, c743_r, c743_a, c743_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I100 (c743_r, c743_a, c743_d, c742_r, c742_a, c742_d, c741_r, c741_a, c741_d);
  BrzSlice_1_34_32 I101 (c740_r, c740_a, c740_d, c739_r, c739_a, c739_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I102 (c739_r, c739_a, c739_d, c738_r, c738_a, c738_d, c737_r, c737_a, c737_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I103 (c736_r, c736_a, c736_d, c735_r, c735_a, c735_d, c733_r, c733_a, c733_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I104 (c735_r, c735_a, c735_d, c734_r, c734_a, c734_d);
  BrzSequence_2_s1_S I105 (c728_r, c728_a, c729_r, c729_a, c730_r, c730_a);
  BrzFetch_33_s5_false I106 (c729_r, c729_a, c726_r, c726_a, c726_d, c731_r, c731_a, c731_d);
  BrzFetch_33_s5_false I107 (c730_r, c730_a, c732_r, c732_a, c732_d, c727_r, c727_a, c727_d);
  BrzVariable_33_1_s0_ I108 (c731_r, c731_a, c731_d, c732_r, c732_a, c732_d);
  BrzCombine_33_32_1 I109 (c726_r, c726_a, c726_d, c725_r, c725_a, c725_d, c721_r, c721_a, c721_d);
  BrzSlice_32_34_1 I110 (c725_r, c725_a, c725_d, c724_r, c724_a, c724_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I111 (c724_r, c724_a, c724_d, c723_r, c723_a, c723_d, c722_r, c722_a, c722_d);
  BrzSlice_1_34_32 I112 (c721_r, c721_a, c721_d, c720_r, c720_a, c720_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I113 (c720_r, c720_a, c720_d, c719_r, c719_a, c719_d, c718_r, c718_a, c718_d);
  BrzSequence_2_s1_S I114 (c713_r, c713_a, c714_r, c714_a, c715_r, c715_a);
  BrzFetch_33_s5_false I115 (c714_r, c714_a, c711_r, c711_a, c711_d, c716_r, c716_a, c716_d);
  BrzFetch_33_s5_false I116 (c715_r, c715_a, c717_r, c717_a, c717_d, c712_r, c712_a, c712_d);
  BrzVariable_33_1_s0_ I117 (c716_r, c716_a, c716_d, c717_r, c717_a, c717_d);
  BrzCombine_33_32_1 I118 (c711_r, c711_a, c711_d, c710_r, c710_a, c710_d, c709_r, c709_a, c709_d);
  BrzCase_1_2_s5_0_3b1 I119 (c704_r, c704_a, c704_d, c659_r, c659_a, c703_r, c703_a);
  BrzFetch_1_s5_false I120 (c705_r, c705_a, c702_r, c702_a, c702_d, c707_r, c707_a, c707_d);
  BrzFetch_1_s5_false I121 (c706_r, c706_a, c708_r, c708_a, c708_d, c704_r, c704_a, c704_d);
  BrzVariable_1_1_s0_ I122 (c707_r, c707_a, c707_d, c708_r, c708_a, c708_d);
  BrzBar_2 I123 (c702_r, c702_a, c702_d, c703_r, c703_a, c682_r, c682_a, c682_d, c701_r, c701_a, c701_d, c674_r, c674_a, c693_r, c693_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I124 (c701_r, c701_a, c701_d, c700_r, c700_a, c700_d, c699_r, c699_a, c699_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I125 (c699_r, c699_a, c699_d, c698_r, c698_a, c698_d);
  BrzSequence_2_s1_S I126 (c693_r, c693_a, c694_r, c694_a, c695_r, c695_a);
  BrzFetch_33_s5_false I127 (c694_r, c694_a, c691_r, c691_a, c691_d, c696_r, c696_a, c696_d);
  BrzFetch_33_s5_false I128 (c695_r, c695_a, c697_r, c697_a, c697_d, c692_r, c692_a, c692_d);
  BrzVariable_33_1_s0_ I129 (c696_r, c696_a, c696_d, c697_r, c697_a, c697_d);
  BrzCombine_33_32_1 I130 (c691_r, c691_a, c691_d, c690_r, c690_a, c690_d, c686_r, c686_a, c686_d);
  BrzSlice_32_34_1 I131 (c690_r, c690_a, c690_d, c689_r, c689_a, c689_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I132 (c689_r, c689_a, c689_d, c688_r, c688_a, c688_d, c687_r, c687_a, c687_d);
  BrzSlice_1_34_32 I133 (c686_r, c686_a, c686_d, c685_r, c685_a, c685_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I134 (c685_r, c685_a, c685_d, c684_r, c684_a, c684_d, c683_r, c683_a, c683_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I135 (c682_r, c682_a, c682_d, c681_r, c681_a, c681_d, c679_r, c679_a, c679_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I136 (c681_r, c681_a, c681_d, c680_r, c680_a, c680_d);
  BrzSequence_2_s1_S I137 (c674_r, c674_a, c675_r, c675_a, c676_r, c676_a);
  BrzFetch_33_s5_false I138 (c675_r, c675_a, c672_r, c672_a, c672_d, c677_r, c677_a, c677_d);
  BrzFetch_33_s5_false I139 (c676_r, c676_a, c678_r, c678_a, c678_d, c673_r, c673_a, c673_d);
  BrzVariable_33_1_s0_ I140 (c677_r, c677_a, c677_d, c678_r, c678_a, c678_d);
  BrzCombine_33_32_1 I141 (c672_r, c672_a, c672_d, c671_r, c671_a, c671_d, c667_r, c667_a, c667_d);
  BrzSlice_32_34_1 I142 (c671_r, c671_a, c671_d, c670_r, c670_a, c670_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I143 (c670_r, c670_a, c670_d, c669_r, c669_a, c669_d, c668_r, c668_a, c668_d);
  BrzSlice_1_34_32 I144 (c667_r, c667_a, c667_d, c666_r, c666_a, c666_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I145 (c666_r, c666_a, c666_d, c665_r, c665_a, c665_d, c664_r, c664_a, c664_d);
  BrzSequence_2_s1_S I146 (c659_r, c659_a, c660_r, c660_a, c661_r, c661_a);
  BrzFetch_33_s5_false I147 (c660_r, c660_a, c657_r, c657_a, c657_d, c662_r, c662_a, c662_d);
  BrzFetch_33_s5_false I148 (c661_r, c661_a, c663_r, c663_a, c663_d, c658_r, c658_a, c658_d);
  BrzVariable_33_1_s0_ I149 (c662_r, c662_a, c662_d, c663_r, c663_a, c663_d);
  BrzCombine_33_32_1 I150 (c657_r, c657_a, c657_d, c656_r, c656_a, c656_d, c655_r, c655_a, c655_d);
  BrzCase_1_2_s5_0_3b1 I151 (c650_r, c650_a, c650_d, c605_r, c605_a, c649_r, c649_a);
  BrzFetch_1_s5_false I152 (c651_r, c651_a, c648_r, c648_a, c648_d, c653_r, c653_a, c653_d);
  BrzFetch_1_s5_false I153 (c652_r, c652_a, c654_r, c654_a, c654_d, c650_r, c650_a, c650_d);
  BrzVariable_1_1_s0_ I154 (c653_r, c653_a, c653_d, c654_r, c654_a, c654_d);
  BrzBar_2 I155 (c648_r, c648_a, c648_d, c649_r, c649_a, c628_r, c628_a, c628_d, c647_r, c647_a, c647_d, c620_r, c620_a, c639_r, c639_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I156 (c647_r, c647_a, c647_d, c646_r, c646_a, c646_d, c645_r, c645_a, c645_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I157 (c645_r, c645_a, c645_d, c644_r, c644_a, c644_d);
  BrzSequence_2_s1_S I158 (c639_r, c639_a, c640_r, c640_a, c641_r, c641_a);
  BrzFetch_33_s5_false I159 (c640_r, c640_a, c637_r, c637_a, c637_d, c642_r, c642_a, c642_d);
  BrzFetch_33_s5_false I160 (c641_r, c641_a, c643_r, c643_a, c643_d, c638_r, c638_a, c638_d);
  BrzVariable_33_1_s0_ I161 (c642_r, c642_a, c642_d, c643_r, c643_a, c643_d);
  BrzCombine_33_32_1 I162 (c637_r, c637_a, c637_d, c636_r, c636_a, c636_d, c632_r, c632_a, c632_d);
  BrzSlice_32_34_1 I163 (c636_r, c636_a, c636_d, c635_r, c635_a, c635_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I164 (c635_r, c635_a, c635_d, c634_r, c634_a, c634_d, c633_r, c633_a, c633_d);
  BrzSlice_1_34_32 I165 (c632_r, c632_a, c632_d, c631_r, c631_a, c631_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I166 (c631_r, c631_a, c631_d, c630_r, c630_a, c630_d, c629_r, c629_a, c629_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I167 (c628_r, c628_a, c628_d, c627_r, c627_a, c627_d, c625_r, c625_a, c625_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I168 (c627_r, c627_a, c627_d, c626_r, c626_a, c626_d);
  BrzSequence_2_s1_S I169 (c620_r, c620_a, c621_r, c621_a, c622_r, c622_a);
  BrzFetch_33_s5_false I170 (c621_r, c621_a, c618_r, c618_a, c618_d, c623_r, c623_a, c623_d);
  BrzFetch_33_s5_false I171 (c622_r, c622_a, c624_r, c624_a, c624_d, c619_r, c619_a, c619_d);
  BrzVariable_33_1_s0_ I172 (c623_r, c623_a, c623_d, c624_r, c624_a, c624_d);
  BrzCombine_33_32_1 I173 (c618_r, c618_a, c618_d, c617_r, c617_a, c617_d, c613_r, c613_a, c613_d);
  BrzSlice_32_34_1 I174 (c617_r, c617_a, c617_d, c616_r, c616_a, c616_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I175 (c616_r, c616_a, c616_d, c615_r, c615_a, c615_d, c614_r, c614_a, c614_d);
  BrzSlice_1_34_32 I176 (c613_r, c613_a, c613_d, c612_r, c612_a, c612_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I177 (c612_r, c612_a, c612_d, c611_r, c611_a, c611_d, c610_r, c610_a, c610_d);
  BrzSequence_2_s1_S I178 (c605_r, c605_a, c606_r, c606_a, c607_r, c607_a);
  BrzFetch_33_s5_false I179 (c606_r, c606_a, c603_r, c603_a, c603_d, c608_r, c608_a, c608_d);
  BrzFetch_33_s5_false I180 (c607_r, c607_a, c609_r, c609_a, c609_d, c604_r, c604_a, c604_d);
  BrzVariable_33_1_s0_ I181 (c608_r, c608_a, c608_d, c609_r, c609_a, c609_d);
  BrzCombine_33_32_1 I182 (c603_r, c603_a, c603_d, c602_r, c602_a, c602_d, c601_r, c601_a, c601_d);
  BrzCase_1_2_s5_0_3b1 I183 (c596_r, c596_a, c596_d, c551_r, c551_a, c595_r, c595_a);
  BrzFetch_1_s5_false I184 (c597_r, c597_a, c594_r, c594_a, c594_d, c599_r, c599_a, c599_d);
  BrzFetch_1_s5_false I185 (c598_r, c598_a, c600_r, c600_a, c600_d, c596_r, c596_a, c596_d);
  BrzVariable_1_1_s0_ I186 (c599_r, c599_a, c599_d, c600_r, c600_a, c600_d);
  BrzBar_2 I187 (c594_r, c594_a, c594_d, c595_r, c595_a, c574_r, c574_a, c574_d, c593_r, c593_a, c593_d, c566_r, c566_a, c585_r, c585_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I188 (c593_r, c593_a, c593_d, c592_r, c592_a, c592_d, c591_r, c591_a, c591_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I189 (c591_r, c591_a, c591_d, c590_r, c590_a, c590_d);
  BrzSequence_2_s1_S I190 (c585_r, c585_a, c586_r, c586_a, c587_r, c587_a);
  BrzFetch_33_s5_false I191 (c586_r, c586_a, c583_r, c583_a, c583_d, c588_r, c588_a, c588_d);
  BrzFetch_33_s5_false I192 (c587_r, c587_a, c589_r, c589_a, c589_d, c584_r, c584_a, c584_d);
  BrzVariable_33_1_s0_ I193 (c588_r, c588_a, c588_d, c589_r, c589_a, c589_d);
  BrzCombine_33_32_1 I194 (c583_r, c583_a, c583_d, c582_r, c582_a, c582_d, c578_r, c578_a, c578_d);
  BrzSlice_32_34_1 I195 (c582_r, c582_a, c582_d, c581_r, c581_a, c581_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I196 (c581_r, c581_a, c581_d, c580_r, c580_a, c580_d, c579_r, c579_a, c579_d);
  BrzSlice_1_34_32 I197 (c578_r, c578_a, c578_d, c577_r, c577_a, c577_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I198 (c577_r, c577_a, c577_d, c576_r, c576_a, c576_d, c575_r, c575_a, c575_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I199 (c574_r, c574_a, c574_d, c573_r, c573_a, c573_d, c571_r, c571_a, c571_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I200 (c573_r, c573_a, c573_d, c572_r, c572_a, c572_d);
  BrzSequence_2_s1_S I201 (c566_r, c566_a, c567_r, c567_a, c568_r, c568_a);
  BrzFetch_33_s5_false I202 (c567_r, c567_a, c564_r, c564_a, c564_d, c569_r, c569_a, c569_d);
  BrzFetch_33_s5_false I203 (c568_r, c568_a, c570_r, c570_a, c570_d, c565_r, c565_a, c565_d);
  BrzVariable_33_1_s0_ I204 (c569_r, c569_a, c569_d, c570_r, c570_a, c570_d);
  BrzCombine_33_32_1 I205 (c564_r, c564_a, c564_d, c563_r, c563_a, c563_d, c559_r, c559_a, c559_d);
  BrzSlice_32_34_1 I206 (c563_r, c563_a, c563_d, c562_r, c562_a, c562_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I207 (c562_r, c562_a, c562_d, c561_r, c561_a, c561_d, c560_r, c560_a, c560_d);
  BrzSlice_1_34_32 I208 (c559_r, c559_a, c559_d, c558_r, c558_a, c558_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I209 (c558_r, c558_a, c558_d, c557_r, c557_a, c557_d, c556_r, c556_a, c556_d);
  BrzSequence_2_s1_S I210 (c551_r, c551_a, c552_r, c552_a, c553_r, c553_a);
  BrzFetch_33_s5_false I211 (c552_r, c552_a, c549_r, c549_a, c549_d, c554_r, c554_a, c554_d);
  BrzFetch_33_s5_false I212 (c553_r, c553_a, c555_r, c555_a, c555_d, c550_r, c550_a, c550_d);
  BrzVariable_33_1_s0_ I213 (c554_r, c554_a, c554_d, c555_r, c555_a, c555_d);
  BrzCombine_33_32_1 I214 (c549_r, c549_a, c549_d, c548_r, c548_a, c548_d, c547_r, c547_a, c547_d);
  BrzCase_1_2_s5_0_3b1 I215 (c542_r, c542_a, c542_d, c497_r, c497_a, c541_r, c541_a);
  BrzFetch_1_s5_false I216 (c543_r, c543_a, c540_r, c540_a, c540_d, c545_r, c545_a, c545_d);
  BrzFetch_1_s5_false I217 (c544_r, c544_a, c546_r, c546_a, c546_d, c542_r, c542_a, c542_d);
  BrzVariable_1_1_s0_ I218 (c545_r, c545_a, c545_d, c546_r, c546_a, c546_d);
  BrzBar_2 I219 (c540_r, c540_a, c540_d, c541_r, c541_a, c520_r, c520_a, c520_d, c539_r, c539_a, c539_d, c512_r, c512_a, c531_r, c531_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I220 (c539_r, c539_a, c539_d, c538_r, c538_a, c538_d, c537_r, c537_a, c537_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I221 (c537_r, c537_a, c537_d, c536_r, c536_a, c536_d);
  BrzSequence_2_s1_S I222 (c531_r, c531_a, c532_r, c532_a, c533_r, c533_a);
  BrzFetch_33_s5_false I223 (c532_r, c532_a, c529_r, c529_a, c529_d, c534_r, c534_a, c534_d);
  BrzFetch_33_s5_false I224 (c533_r, c533_a, c535_r, c535_a, c535_d, c530_r, c530_a, c530_d);
  BrzVariable_33_1_s0_ I225 (c534_r, c534_a, c534_d, c535_r, c535_a, c535_d);
  BrzCombine_33_32_1 I226 (c529_r, c529_a, c529_d, c528_r, c528_a, c528_d, c524_r, c524_a, c524_d);
  BrzSlice_32_34_1 I227 (c528_r, c528_a, c528_d, c527_r, c527_a, c527_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I228 (c527_r, c527_a, c527_d, c526_r, c526_a, c526_d, c525_r, c525_a, c525_d);
  BrzSlice_1_34_32 I229 (c524_r, c524_a, c524_d, c523_r, c523_a, c523_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I230 (c523_r, c523_a, c523_d, c522_r, c522_a, c522_d, c521_r, c521_a, c521_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I231 (c520_r, c520_a, c520_d, c519_r, c519_a, c519_d, c517_r, c517_a, c517_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I232 (c519_r, c519_a, c519_d, c518_r, c518_a, c518_d);
  BrzSequence_2_s1_S I233 (c512_r, c512_a, c513_r, c513_a, c514_r, c514_a);
  BrzFetch_33_s5_false I234 (c513_r, c513_a, c510_r, c510_a, c510_d, c515_r, c515_a, c515_d);
  BrzFetch_33_s5_false I235 (c514_r, c514_a, c516_r, c516_a, c516_d, c511_r, c511_a, c511_d);
  BrzVariable_33_1_s0_ I236 (c515_r, c515_a, c515_d, c516_r, c516_a, c516_d);
  BrzCombine_33_32_1 I237 (c510_r, c510_a, c510_d, c509_r, c509_a, c509_d, c505_r, c505_a, c505_d);
  BrzSlice_32_34_1 I238 (c509_r, c509_a, c509_d, c508_r, c508_a, c508_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I239 (c508_r, c508_a, c508_d, c507_r, c507_a, c507_d, c506_r, c506_a, c506_d);
  BrzSlice_1_34_32 I240 (c505_r, c505_a, c505_d, c504_r, c504_a, c504_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I241 (c504_r, c504_a, c504_d, c503_r, c503_a, c503_d, c502_r, c502_a, c502_d);
  BrzSequence_2_s1_S I242 (c497_r, c497_a, c498_r, c498_a, c499_r, c499_a);
  BrzFetch_33_s5_false I243 (c498_r, c498_a, c495_r, c495_a, c495_d, c500_r, c500_a, c500_d);
  BrzFetch_33_s5_false I244 (c499_r, c499_a, c501_r, c501_a, c501_d, c496_r, c496_a, c496_d);
  BrzVariable_33_1_s0_ I245 (c500_r, c500_a, c500_d, c501_r, c501_a, c501_d);
  BrzCombine_33_32_1 I246 (c495_r, c495_a, c495_d, c494_r, c494_a, c494_d, c493_r, c493_a, c493_d);
  BrzCase_1_2_s5_0_3b1 I247 (c488_r, c488_a, c488_d, c443_r, c443_a, c487_r, c487_a);
  BrzFetch_1_s5_false I248 (c489_r, c489_a, c486_r, c486_a, c486_d, c491_r, c491_a, c491_d);
  BrzFetch_1_s5_false I249 (c490_r, c490_a, c492_r, c492_a, c492_d, c488_r, c488_a, c488_d);
  BrzVariable_1_1_s0_ I250 (c491_r, c491_a, c491_d, c492_r, c492_a, c492_d);
  BrzBar_2 I251 (c486_r, c486_a, c486_d, c487_r, c487_a, c466_r, c466_a, c466_d, c485_r, c485_a, c485_d, c458_r, c458_a, c477_r, c477_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I252 (c485_r, c485_a, c485_d, c484_r, c484_a, c484_d, c483_r, c483_a, c483_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I253 (c483_r, c483_a, c483_d, c482_r, c482_a, c482_d);
  BrzSequence_2_s1_S I254 (c477_r, c477_a, c478_r, c478_a, c479_r, c479_a);
  BrzFetch_33_s5_false I255 (c478_r, c478_a, c475_r, c475_a, c475_d, c480_r, c480_a, c480_d);
  BrzFetch_33_s5_false I256 (c479_r, c479_a, c481_r, c481_a, c481_d, c476_r, c476_a, c476_d);
  BrzVariable_33_1_s0_ I257 (c480_r, c480_a, c480_d, c481_r, c481_a, c481_d);
  BrzCombine_33_32_1 I258 (c475_r, c475_a, c475_d, c474_r, c474_a, c474_d, c470_r, c470_a, c470_d);
  BrzSlice_32_34_1 I259 (c474_r, c474_a, c474_d, c473_r, c473_a, c473_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I260 (c473_r, c473_a, c473_d, c472_r, c472_a, c472_d, c471_r, c471_a, c471_d);
  BrzSlice_1_34_32 I261 (c470_r, c470_a, c470_d, c469_r, c469_a, c469_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I262 (c469_r, c469_a, c469_d, c468_r, c468_a, c468_d, c467_r, c467_a, c467_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I263 (c466_r, c466_a, c466_d, c465_r, c465_a, c465_d, c463_r, c463_a, c463_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I264 (c465_r, c465_a, c465_d, c464_r, c464_a, c464_d);
  BrzSequence_2_s1_S I265 (c458_r, c458_a, c459_r, c459_a, c460_r, c460_a);
  BrzFetch_33_s5_false I266 (c459_r, c459_a, c456_r, c456_a, c456_d, c461_r, c461_a, c461_d);
  BrzFetch_33_s5_false I267 (c460_r, c460_a, c462_r, c462_a, c462_d, c457_r, c457_a, c457_d);
  BrzVariable_33_1_s0_ I268 (c461_r, c461_a, c461_d, c462_r, c462_a, c462_d);
  BrzCombine_33_32_1 I269 (c456_r, c456_a, c456_d, c455_r, c455_a, c455_d, c451_r, c451_a, c451_d);
  BrzSlice_32_34_1 I270 (c455_r, c455_a, c455_d, c454_r, c454_a, c454_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I271 (c454_r, c454_a, c454_d, c453_r, c453_a, c453_d, c452_r, c452_a, c452_d);
  BrzSlice_1_34_32 I272 (c451_r, c451_a, c451_d, c450_r, c450_a, c450_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I273 (c450_r, c450_a, c450_d, c449_r, c449_a, c449_d, c448_r, c448_a, c448_d);
  BrzSequence_2_s1_S I274 (c443_r, c443_a, c444_r, c444_a, c445_r, c445_a);
  BrzFetch_33_s5_false I275 (c444_r, c444_a, c441_r, c441_a, c441_d, c446_r, c446_a, c446_d);
  BrzFetch_33_s5_false I276 (c445_r, c445_a, c447_r, c447_a, c447_d, c442_r, c442_a, c442_d);
  BrzVariable_33_1_s0_ I277 (c446_r, c446_a, c446_d, c447_r, c447_a, c447_d);
  BrzCombine_33_32_1 I278 (c441_r, c441_a, c441_d, c440_r, c440_a, c440_d, c439_r, c439_a, c439_d);
  BrzCase_1_2_s5_0_3b1 I279 (c434_r, c434_a, c434_d, c389_r, c389_a, c433_r, c433_a);
  BrzFetch_1_s5_false I280 (c435_r, c435_a, c432_r, c432_a, c432_d, c437_r, c437_a, c437_d);
  BrzFetch_1_s5_false I281 (c436_r, c436_a, c438_r, c438_a, c438_d, c434_r, c434_a, c434_d);
  BrzVariable_1_1_s0_ I282 (c437_r, c437_a, c437_d, c438_r, c438_a, c438_d);
  BrzBar_2 I283 (c432_r, c432_a, c432_d, c433_r, c433_a, c412_r, c412_a, c412_d, c431_r, c431_a, c431_d, c404_r, c404_a, c423_r, c423_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I284 (c431_r, c431_a, c431_d, c430_r, c430_a, c430_d, c429_r, c429_a, c429_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I285 (c429_r, c429_a, c429_d, c428_r, c428_a, c428_d);
  BrzSequence_2_s1_S I286 (c423_r, c423_a, c424_r, c424_a, c425_r, c425_a);
  BrzFetch_33_s5_false I287 (c424_r, c424_a, c421_r, c421_a, c421_d, c426_r, c426_a, c426_d);
  BrzFetch_33_s5_false I288 (c425_r, c425_a, c427_r, c427_a, c427_d, c422_r, c422_a, c422_d);
  BrzVariable_33_1_s0_ I289 (c426_r, c426_a, c426_d, c427_r, c427_a, c427_d);
  BrzCombine_33_32_1 I290 (c421_r, c421_a, c421_d, c420_r, c420_a, c420_d, c416_r, c416_a, c416_d);
  BrzSlice_32_34_1 I291 (c420_r, c420_a, c420_d, c419_r, c419_a, c419_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I292 (c419_r, c419_a, c419_d, c418_r, c418_a, c418_d, c417_r, c417_a, c417_d);
  BrzSlice_1_34_32 I293 (c416_r, c416_a, c416_d, c415_r, c415_a, c415_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I294 (c415_r, c415_a, c415_d, c414_r, c414_a, c414_d, c413_r, c413_a, c413_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I295 (c412_r, c412_a, c412_d, c411_r, c411_a, c411_d, c409_r, c409_a, c409_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I296 (c411_r, c411_a, c411_d, c410_r, c410_a, c410_d);
  BrzSequence_2_s1_S I297 (c404_r, c404_a, c405_r, c405_a, c406_r, c406_a);
  BrzFetch_33_s5_false I298 (c405_r, c405_a, c402_r, c402_a, c402_d, c407_r, c407_a, c407_d);
  BrzFetch_33_s5_false I299 (c406_r, c406_a, c408_r, c408_a, c408_d, c403_r, c403_a, c403_d);
  BrzVariable_33_1_s0_ I300 (c407_r, c407_a, c407_d, c408_r, c408_a, c408_d);
  BrzCombine_33_32_1 I301 (c402_r, c402_a, c402_d, c401_r, c401_a, c401_d, c397_r, c397_a, c397_d);
  BrzSlice_32_34_1 I302 (c401_r, c401_a, c401_d, c400_r, c400_a, c400_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I303 (c400_r, c400_a, c400_d, c399_r, c399_a, c399_d, c398_r, c398_a, c398_d);
  BrzSlice_1_34_32 I304 (c397_r, c397_a, c397_d, c396_r, c396_a, c396_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I305 (c396_r, c396_a, c396_d, c395_r, c395_a, c395_d, c394_r, c394_a, c394_d);
  BrzSequence_2_s1_S I306 (c389_r, c389_a, c390_r, c390_a, c391_r, c391_a);
  BrzFetch_33_s5_false I307 (c390_r, c390_a, c387_r, c387_a, c387_d, c392_r, c392_a, c392_d);
  BrzFetch_33_s5_false I308 (c391_r, c391_a, c393_r, c393_a, c393_d, c388_r, c388_a, c388_d);
  BrzVariable_33_1_s0_ I309 (c392_r, c392_a, c392_d, c393_r, c393_a, c393_d);
  BrzCombine_33_32_1 I310 (c387_r, c387_a, c387_d, c386_r, c386_a, c386_d, c385_r, c385_a, c385_d);
  BrzCase_1_2_s5_0_3b1 I311 (c380_r, c380_a, c380_d, c335_r, c335_a, c379_r, c379_a);
  BrzFetch_1_s5_false I312 (c381_r, c381_a, c378_r, c378_a, c378_d, c383_r, c383_a, c383_d);
  BrzFetch_1_s5_false I313 (c382_r, c382_a, c384_r, c384_a, c384_d, c380_r, c380_a, c380_d);
  BrzVariable_1_1_s0_ I314 (c383_r, c383_a, c383_d, c384_r, c384_a, c384_d);
  BrzBar_2 I315 (c378_r, c378_a, c378_d, c379_r, c379_a, c358_r, c358_a, c358_d, c377_r, c377_a, c377_d, c350_r, c350_a, c369_r, c369_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I316 (c377_r, c377_a, c377_d, c376_r, c376_a, c376_d, c375_r, c375_a, c375_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I317 (c375_r, c375_a, c375_d, c374_r, c374_a, c374_d);
  BrzSequence_2_s1_S I318 (c369_r, c369_a, c370_r, c370_a, c371_r, c371_a);
  BrzFetch_33_s5_false I319 (c370_r, c370_a, c367_r, c367_a, c367_d, c372_r, c372_a, c372_d);
  BrzFetch_33_s5_false I320 (c371_r, c371_a, c373_r, c373_a, c373_d, c368_r, c368_a, c368_d);
  BrzVariable_33_1_s0_ I321 (c372_r, c372_a, c372_d, c373_r, c373_a, c373_d);
  BrzCombine_33_32_1 I322 (c367_r, c367_a, c367_d, c366_r, c366_a, c366_d, c362_r, c362_a, c362_d);
  BrzSlice_32_34_1 I323 (c366_r, c366_a, c366_d, c365_r, c365_a, c365_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I324 (c365_r, c365_a, c365_d, c364_r, c364_a, c364_d, c363_r, c363_a, c363_d);
  BrzSlice_1_34_32 I325 (c362_r, c362_a, c362_d, c361_r, c361_a, c361_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I326 (c361_r, c361_a, c361_d, c360_r, c360_a, c360_d, c359_r, c359_a, c359_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I327 (c358_r, c358_a, c358_d, c357_r, c357_a, c357_d, c355_r, c355_a, c355_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I328 (c357_r, c357_a, c357_d, c356_r, c356_a, c356_d);
  BrzSequence_2_s1_S I329 (c350_r, c350_a, c351_r, c351_a, c352_r, c352_a);
  BrzFetch_33_s5_false I330 (c351_r, c351_a, c348_r, c348_a, c348_d, c353_r, c353_a, c353_d);
  BrzFetch_33_s5_false I331 (c352_r, c352_a, c354_r, c354_a, c354_d, c349_r, c349_a, c349_d);
  BrzVariable_33_1_s0_ I332 (c353_r, c353_a, c353_d, c354_r, c354_a, c354_d);
  BrzCombine_33_32_1 I333 (c348_r, c348_a, c348_d, c347_r, c347_a, c347_d, c343_r, c343_a, c343_d);
  BrzSlice_32_34_1 I334 (c347_r, c347_a, c347_d, c346_r, c346_a, c346_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I335 (c346_r, c346_a, c346_d, c345_r, c345_a, c345_d, c344_r, c344_a, c344_d);
  BrzSlice_1_34_32 I336 (c343_r, c343_a, c343_d, c342_r, c342_a, c342_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I337 (c342_r, c342_a, c342_d, c341_r, c341_a, c341_d, c340_r, c340_a, c340_d);
  BrzSequence_2_s1_S I338 (c335_r, c335_a, c336_r, c336_a, c337_r, c337_a);
  BrzFetch_33_s5_false I339 (c336_r, c336_a, c333_r, c333_a, c333_d, c338_r, c338_a, c338_d);
  BrzFetch_33_s5_false I340 (c337_r, c337_a, c339_r, c339_a, c339_d, c334_r, c334_a, c334_d);
  BrzVariable_33_1_s0_ I341 (c338_r, c338_a, c338_d, c339_r, c339_a, c339_d);
  BrzCombine_33_32_1 I342 (c333_r, c333_a, c333_d, c332_r, c332_a, c332_d, c331_r, c331_a, c331_d);
  BrzCase_1_2_s5_0_3b1 I343 (c326_r, c326_a, c326_d, c281_r, c281_a, c325_r, c325_a);
  BrzFetch_1_s5_false I344 (c327_r, c327_a, c324_r, c324_a, c324_d, c329_r, c329_a, c329_d);
  BrzFetch_1_s5_false I345 (c328_r, c328_a, c330_r, c330_a, c330_d, c326_r, c326_a, c326_d);
  BrzVariable_1_1_s0_ I346 (c329_r, c329_a, c329_d, c330_r, c330_a, c330_d);
  BrzBar_2 I347 (c324_r, c324_a, c324_d, c325_r, c325_a, c304_r, c304_a, c304_d, c323_r, c323_a, c323_d, c296_r, c296_a, c315_r, c315_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I348 (c323_r, c323_a, c323_d, c322_r, c322_a, c322_d, c321_r, c321_a, c321_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I349 (c321_r, c321_a, c321_d, c320_r, c320_a, c320_d);
  BrzSequence_2_s1_S I350 (c315_r, c315_a, c316_r, c316_a, c317_r, c317_a);
  BrzFetch_33_s5_false I351 (c316_r, c316_a, c313_r, c313_a, c313_d, c318_r, c318_a, c318_d);
  BrzFetch_33_s5_false I352 (c317_r, c317_a, c319_r, c319_a, c319_d, c314_r, c314_a, c314_d);
  BrzVariable_33_1_s0_ I353 (c318_r, c318_a, c318_d, c319_r, c319_a, c319_d);
  BrzCombine_33_32_1 I354 (c313_r, c313_a, c313_d, c312_r, c312_a, c312_d, c308_r, c308_a, c308_d);
  BrzSlice_32_34_1 I355 (c312_r, c312_a, c312_d, c311_r, c311_a, c311_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I356 (c311_r, c311_a, c311_d, c310_r, c310_a, c310_d, c309_r, c309_a, c309_d);
  BrzSlice_1_34_32 I357 (c308_r, c308_a, c308_d, c307_r, c307_a, c307_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I358 (c307_r, c307_a, c307_d, c306_r, c306_a, c306_d, c305_r, c305_a, c305_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I359 (c304_r, c304_a, c304_d, c303_r, c303_a, c303_d, c301_r, c301_a, c301_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I360 (c303_r, c303_a, c303_d, c302_r, c302_a, c302_d);
  BrzSequence_2_s1_S I361 (c296_r, c296_a, c297_r, c297_a, c298_r, c298_a);
  BrzFetch_33_s5_false I362 (c297_r, c297_a, c294_r, c294_a, c294_d, c299_r, c299_a, c299_d);
  BrzFetch_33_s5_false I363 (c298_r, c298_a, c300_r, c300_a, c300_d, c295_r, c295_a, c295_d);
  BrzVariable_33_1_s0_ I364 (c299_r, c299_a, c299_d, c300_r, c300_a, c300_d);
  BrzCombine_33_32_1 I365 (c294_r, c294_a, c294_d, c293_r, c293_a, c293_d, c289_r, c289_a, c289_d);
  BrzSlice_32_34_1 I366 (c293_r, c293_a, c293_d, c292_r, c292_a, c292_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I367 (c292_r, c292_a, c292_d, c291_r, c291_a, c291_d, c290_r, c290_a, c290_d);
  BrzSlice_1_34_32 I368 (c289_r, c289_a, c289_d, c288_r, c288_a, c288_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I369 (c288_r, c288_a, c288_d, c287_r, c287_a, c287_d, c286_r, c286_a, c286_d);
  BrzSequence_2_s1_S I370 (c281_r, c281_a, c282_r, c282_a, c283_r, c283_a);
  BrzFetch_33_s5_false I371 (c282_r, c282_a, c279_r, c279_a, c279_d, c284_r, c284_a, c284_d);
  BrzFetch_33_s5_false I372 (c283_r, c283_a, c285_r, c285_a, c285_d, c280_r, c280_a, c280_d);
  BrzVariable_33_1_s0_ I373 (c284_r, c284_a, c284_d, c285_r, c285_a, c285_d);
  BrzCombine_33_32_1 I374 (c279_r, c279_a, c279_d, c278_r, c278_a, c278_d, c277_r, c277_a, c277_d);
  BrzCase_1_2_s5_0_3b1 I375 (c272_r, c272_a, c272_d, c227_r, c227_a, c271_r, c271_a);
  BrzFetch_1_s5_false I376 (c273_r, c273_a, c270_r, c270_a, c270_d, c275_r, c275_a, c275_d);
  BrzFetch_1_s5_false I377 (c274_r, c274_a, c276_r, c276_a, c276_d, c272_r, c272_a, c272_d);
  BrzVariable_1_1_s0_ I378 (c275_r, c275_a, c275_d, c276_r, c276_a, c276_d);
  BrzBar_2 I379 (c270_r, c270_a, c270_d, c271_r, c271_a, c250_r, c250_a, c250_d, c269_r, c269_a, c269_d, c242_r, c242_a, c261_r, c261_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I380 (c269_r, c269_a, c269_d, c268_r, c268_a, c268_d, c267_r, c267_a, c267_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I381 (c267_r, c267_a, c267_d, c266_r, c266_a, c266_d);
  BrzSequence_2_s1_S I382 (c261_r, c261_a, c262_r, c262_a, c263_r, c263_a);
  BrzFetch_33_s5_false I383 (c262_r, c262_a, c259_r, c259_a, c259_d, c264_r, c264_a, c264_d);
  BrzFetch_33_s5_false I384 (c263_r, c263_a, c265_r, c265_a, c265_d, c260_r, c260_a, c260_d);
  BrzVariable_33_1_s0_ I385 (c264_r, c264_a, c264_d, c265_r, c265_a, c265_d);
  BrzCombine_33_32_1 I386 (c259_r, c259_a, c259_d, c258_r, c258_a, c258_d, c254_r, c254_a, c254_d);
  BrzSlice_32_34_1 I387 (c258_r, c258_a, c258_d, c257_r, c257_a, c257_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I388 (c257_r, c257_a, c257_d, c256_r, c256_a, c256_d, c255_r, c255_a, c255_d);
  BrzSlice_1_34_32 I389 (c254_r, c254_a, c254_d, c253_r, c253_a, c253_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I390 (c253_r, c253_a, c253_d, c252_r, c252_a, c252_d, c251_r, c251_a, c251_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I391 (c250_r, c250_a, c250_d, c249_r, c249_a, c249_d, c247_r, c247_a, c247_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I392 (c249_r, c249_a, c249_d, c248_r, c248_a, c248_d);
  BrzSequence_2_s1_S I393 (c242_r, c242_a, c243_r, c243_a, c244_r, c244_a);
  BrzFetch_33_s5_false I394 (c243_r, c243_a, c240_r, c240_a, c240_d, c245_r, c245_a, c245_d);
  BrzFetch_33_s5_false I395 (c244_r, c244_a, c246_r, c246_a, c246_d, c241_r, c241_a, c241_d);
  BrzVariable_33_1_s0_ I396 (c245_r, c245_a, c245_d, c246_r, c246_a, c246_d);
  BrzCombine_33_32_1 I397 (c240_r, c240_a, c240_d, c239_r, c239_a, c239_d, c235_r, c235_a, c235_d);
  BrzSlice_32_34_1 I398 (c239_r, c239_a, c239_d, c238_r, c238_a, c238_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I399 (c238_r, c238_a, c238_d, c237_r, c237_a, c237_d, c236_r, c236_a, c236_d);
  BrzSlice_1_34_32 I400 (c235_r, c235_a, c235_d, c234_r, c234_a, c234_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I401 (c234_r, c234_a, c234_d, c233_r, c233_a, c233_d, c232_r, c232_a, c232_d);
  BrzSequence_2_s1_S I402 (c227_r, c227_a, c228_r, c228_a, c229_r, c229_a);
  BrzFetch_33_s5_false I403 (c228_r, c228_a, c225_r, c225_a, c225_d, c230_r, c230_a, c230_d);
  BrzFetch_33_s5_false I404 (c229_r, c229_a, c231_r, c231_a, c231_d, c226_r, c226_a, c226_d);
  BrzVariable_33_1_s0_ I405 (c230_r, c230_a, c230_d, c231_r, c231_a, c231_d);
  BrzCombine_33_32_1 I406 (c225_r, c225_a, c225_d, c224_r, c224_a, c224_d, c223_r, c223_a, c223_d);
  BrzCase_1_2_s5_0_3b1 I407 (c218_r, c218_a, c218_d, c173_r, c173_a, c217_r, c217_a);
  BrzFetch_1_s5_false I408 (c219_r, c219_a, c216_r, c216_a, c216_d, c221_r, c221_a, c221_d);
  BrzFetch_1_s5_false I409 (c220_r, c220_a, c222_r, c222_a, c222_d, c218_r, c218_a, c218_d);
  BrzVariable_1_1_s0_ I410 (c221_r, c221_a, c221_d, c222_r, c222_a, c222_d);
  BrzBar_2 I411 (c216_r, c216_a, c216_d, c217_r, c217_a, c196_r, c196_a, c196_d, c215_r, c215_a, c215_d, c188_r, c188_a, c207_r, c207_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I412 (c215_r, c215_a, c215_d, c214_r, c214_a, c214_d, c213_r, c213_a, c213_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I413 (c213_r, c213_a, c213_d, c212_r, c212_a, c212_d);
  BrzSequence_2_s1_S I414 (c207_r, c207_a, c208_r, c208_a, c209_r, c209_a);
  BrzFetch_33_s5_false I415 (c208_r, c208_a, c205_r, c205_a, c205_d, c210_r, c210_a, c210_d);
  BrzFetch_33_s5_false I416 (c209_r, c209_a, c211_r, c211_a, c211_d, c206_r, c206_a, c206_d);
  BrzVariable_33_1_s0_ I417 (c210_r, c210_a, c210_d, c211_r, c211_a, c211_d);
  BrzCombine_33_32_1 I418 (c205_r, c205_a, c205_d, c204_r, c204_a, c204_d, c200_r, c200_a, c200_d);
  BrzSlice_32_34_1 I419 (c204_r, c204_a, c204_d, c203_r, c203_a, c203_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I420 (c203_r, c203_a, c203_d, c202_r, c202_a, c202_d, c201_r, c201_a, c201_d);
  BrzSlice_1_34_32 I421 (c200_r, c200_a, c200_d, c199_r, c199_a, c199_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I422 (c199_r, c199_a, c199_d, c198_r, c198_a, c198_d, c197_r, c197_a, c197_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I423 (c196_r, c196_a, c196_d, c195_r, c195_a, c195_d, c193_r, c193_a, c193_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I424 (c195_r, c195_a, c195_d, c194_r, c194_a, c194_d);
  BrzSequence_2_s1_S I425 (c188_r, c188_a, c189_r, c189_a, c190_r, c190_a);
  BrzFetch_33_s5_false I426 (c189_r, c189_a, c186_r, c186_a, c186_d, c191_r, c191_a, c191_d);
  BrzFetch_33_s5_false I427 (c190_r, c190_a, c192_r, c192_a, c192_d, c187_r, c187_a, c187_d);
  BrzVariable_33_1_s0_ I428 (c191_r, c191_a, c191_d, c192_r, c192_a, c192_d);
  BrzCombine_33_32_1 I429 (c186_r, c186_a, c186_d, c185_r, c185_a, c185_d, c181_r, c181_a, c181_d);
  BrzSlice_32_34_1 I430 (c185_r, c185_a, c185_d, c184_r, c184_a, c184_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I431 (c184_r, c184_a, c184_d, c183_r, c183_a, c183_d, c182_r, c182_a, c182_d);
  BrzSlice_1_34_32 I432 (c181_r, c181_a, c181_d, c180_r, c180_a, c180_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I433 (c180_r, c180_a, c180_d, c179_r, c179_a, c179_d, c178_r, c178_a, c178_d);
  BrzSequence_2_s1_S I434 (c173_r, c173_a, c174_r, c174_a, c175_r, c175_a);
  BrzFetch_33_s5_false I435 (c174_r, c174_a, c171_r, c171_a, c171_d, c176_r, c176_a, c176_d);
  BrzFetch_33_s5_false I436 (c175_r, c175_a, c177_r, c177_a, c177_d, c172_r, c172_a, c172_d);
  BrzVariable_33_1_s0_ I437 (c176_r, c176_a, c176_d, c177_r, c177_a, c177_d);
  BrzCombine_33_32_1 I438 (c171_r, c171_a, c171_d, c170_r, c170_a, c170_d, c169_r, c169_a, c169_d);
  BrzCase_1_2_s5_0_3b1 I439 (c164_r, c164_a, c164_d, c119_r, c119_a, c163_r, c163_a);
  BrzFetch_1_s5_false I440 (c165_r, c165_a, c162_r, c162_a, c162_d, c167_r, c167_a, c167_d);
  BrzFetch_1_s5_false I441 (c166_r, c166_a, c168_r, c168_a, c168_d, c164_r, c164_a, c164_d);
  BrzVariable_1_1_s0_ I442 (c167_r, c167_a, c167_d, c168_r, c168_a, c168_d);
  BrzBar_2 I443 (c162_r, c162_a, c162_d, c163_r, c163_a, c142_r, c142_a, c142_d, c161_r, c161_a, c161_d, c134_r, c134_a, c153_r, c153_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I444 (c161_r, c161_a, c161_d, c160_r, c160_a, c160_d, c159_r, c159_a, c159_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I445 (c159_r, c159_a, c159_d, c158_r, c158_a, c158_d);
  BrzSequence_2_s1_S I446 (c153_r, c153_a, c154_r, c154_a, c155_r, c155_a);
  BrzFetch_33_s5_false I447 (c154_r, c154_a, c151_r, c151_a, c151_d, c156_r, c156_a, c156_d);
  BrzFetch_33_s5_false I448 (c155_r, c155_a, c157_r, c157_a, c157_d, c152_r, c152_a, c152_d);
  BrzVariable_33_1_s0_ I449 (c156_r, c156_a, c156_d, c157_r, c157_a, c157_d);
  BrzCombine_33_32_1 I450 (c151_r, c151_a, c151_d, c150_r, c150_a, c150_d, c146_r, c146_a, c146_d);
  BrzSlice_32_34_1 I451 (c150_r, c150_a, c150_d, c149_r, c149_a, c149_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I452 (c149_r, c149_a, c149_d, c148_r, c148_a, c148_d, c147_r, c147_a, c147_d);
  BrzSlice_1_34_32 I453 (c146_r, c146_a, c146_d, c145_r, c145_a, c145_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I454 (c145_r, c145_a, c145_d, c144_r, c144_a, c144_d, c143_r, c143_a, c143_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I455 (c142_r, c142_a, c142_d, c141_r, c141_a, c141_d, c139_r, c139_a, c139_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I456 (c141_r, c141_a, c141_d, c140_r, c140_a, c140_d);
  BrzSequence_2_s1_S I457 (c134_r, c134_a, c135_r, c135_a, c136_r, c136_a);
  BrzFetch_33_s5_false I458 (c135_r, c135_a, c132_r, c132_a, c132_d, c137_r, c137_a, c137_d);
  BrzFetch_33_s5_false I459 (c136_r, c136_a, c138_r, c138_a, c138_d, c133_r, c133_a, c133_d);
  BrzVariable_33_1_s0_ I460 (c137_r, c137_a, c137_d, c138_r, c138_a, c138_d);
  BrzCombine_33_32_1 I461 (c132_r, c132_a, c132_d, c131_r, c131_a, c131_d, c127_r, c127_a, c127_d);
  BrzSlice_32_34_1 I462 (c131_r, c131_a, c131_d, c130_r, c130_a, c130_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I463 (c130_r, c130_a, c130_d, c129_r, c129_a, c129_d, c128_r, c128_a, c128_d);
  BrzSlice_1_34_32 I464 (c127_r, c127_a, c127_d, c126_r, c126_a, c126_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I465 (c126_r, c126_a, c126_d, c125_r, c125_a, c125_d, c124_r, c124_a, c124_d);
  BrzSequence_2_s1_S I466 (c119_r, c119_a, c120_r, c120_a, c121_r, c121_a);
  BrzFetch_33_s5_false I467 (c120_r, c120_a, c117_r, c117_a, c117_d, c122_r, c122_a, c122_d);
  BrzFetch_33_s5_false I468 (c121_r, c121_a, c123_r, c123_a, c123_d, c118_r, c118_a, c118_d);
  BrzVariable_33_1_s0_ I469 (c122_r, c122_a, c122_d, c123_r, c123_a, c123_d);
  BrzCombine_33_32_1 I470 (c117_r, c117_a, c117_d, c116_r, c116_a, c116_d, c115_r, c115_a, c115_d);
  BrzCase_1_2_s5_0_3b1 I471 (c110_r, c110_a, c110_d, c65_r, c65_a, c109_r, c109_a);
  BrzFetch_1_s5_false I472 (c111_r, c111_a, c108_r, c108_a, c108_d, c113_r, c113_a, c113_d);
  BrzFetch_1_s5_false I473 (c112_r, c112_a, c114_r, c114_a, c114_d, c110_r, c110_a, c110_d);
  BrzVariable_1_1_s0_ I474 (c113_r, c113_a, c113_d, c114_r, c114_a, c114_d);
  BrzBar_2 I475 (c108_r, c108_a, c108_d, c109_r, c109_a, c88_r, c88_a, c88_d, c107_r, c107_a, c107_d, c80_r, c80_a, c99_r, c99_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I476 (c107_r, c107_a, c107_d, c106_r, c106_a, c106_d, c105_r, c105_a, c105_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I477 (c105_r, c105_a, c105_d, c104_r, c104_a, c104_d);
  BrzSequence_2_s1_S I478 (c99_r, c99_a, c100_r, c100_a, c101_r, c101_a);
  BrzFetch_33_s5_false I479 (c100_r, c100_a, c97_r, c97_a, c97_d, c102_r, c102_a, c102_d);
  BrzFetch_33_s5_false I480 (c101_r, c101_a, c103_r, c103_a, c103_d, c98_r, c98_a, c98_d);
  BrzVariable_33_1_s0_ I481 (c102_r, c102_a, c102_d, c103_r, c103_a, c103_d);
  BrzCombine_33_32_1 I482 (c97_r, c97_a, c97_d, c96_r, c96_a, c96_d, c92_r, c92_a, c92_d);
  BrzSlice_32_34_1 I483 (c96_r, c96_a, c96_d, c95_r, c95_a, c95_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I484 (c95_r, c95_a, c95_d, c94_r, c94_a, c94_d, c93_r, c93_a, c93_d);
  BrzSlice_1_34_32 I485 (c92_r, c92_a, c92_d, c91_r, c91_a, c91_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I486 (c91_r, c91_a, c91_d, c90_r, c90_a, c90_d, c89_r, c89_a, c89_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I487 (c88_r, c88_a, c88_d, c87_r, c87_a, c87_d, c85_r, c85_a, c85_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I488 (c87_r, c87_a, c87_d, c86_r, c86_a, c86_d);
  BrzSequence_2_s1_S I489 (c80_r, c80_a, c81_r, c81_a, c82_r, c82_a);
  BrzFetch_33_s5_false I490 (c81_r, c81_a, c78_r, c78_a, c78_d, c83_r, c83_a, c83_d);
  BrzFetch_33_s5_false I491 (c82_r, c82_a, c84_r, c84_a, c84_d, c79_r, c79_a, c79_d);
  BrzVariable_33_1_s0_ I492 (c83_r, c83_a, c83_d, c84_r, c84_a, c84_d);
  BrzCombine_33_32_1 I493 (c78_r, c78_a, c78_d, c77_r, c77_a, c77_d, c73_r, c73_a, c73_d);
  BrzSlice_32_34_1 I494 (c77_r, c77_a, c77_d, c76_r, c76_a, c76_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I495 (c76_r, c76_a, c76_d, c75_r, c75_a, c75_d, c74_r, c74_a, c74_d);
  BrzSlice_1_34_32 I496 (c73_r, c73_a, c73_d, c72_r, c72_a, c72_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I497 (c72_r, c72_a, c72_d, c71_r, c71_a, c71_d, c70_r, c70_a, c70_d);
  BrzSequence_2_s1_S I498 (c65_r, c65_a, c66_r, c66_a, c67_r, c67_a);
  BrzFetch_33_s5_false I499 (c66_r, c66_a, c63_r, c63_a, c63_d, c68_r, c68_a, c68_d);
  BrzFetch_33_s5_false I500 (c67_r, c67_a, c69_r, c69_a, c69_d, c64_r, c64_a, c64_d);
  BrzVariable_33_1_s0_ I501 (c68_r, c68_a, c68_d, c69_r, c69_a, c69_d);
  BrzCombine_33_32_1 I502 (c63_r, c63_a, c63_d, c62_r, c62_a, c62_d, c61_r, c61_a, c61_d);
  BrzCase_1_2_s5_0_3b1 I503 (c56_r, c56_a, c56_d, c11_r, c11_a, c55_r, c55_a);
  BrzFetch_1_s5_false I504 (c57_r, c57_a, c54_r, c54_a, c54_d, c59_r, c59_a, c59_d);
  BrzFetch_1_s5_false I505 (c58_r, c58_a, c60_r, c60_a, c60_d, c56_r, c56_a, c56_d);
  BrzVariable_1_1_s0_ I506 (c59_r, c59_a, c59_d, c60_r, c60_a, c60_d);
  BrzBar_2 I507 (c54_r, c54_a, c54_d, c55_r, c55_a, c34_r, c34_a, c34_d, c53_r, c53_a, c53_d, c26_r, c26_a, c45_r, c45_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I508 (c53_r, c53_a, c53_d, c52_r, c52_a, c52_d, c51_r, c51_a, c51_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I509 (c51_r, c51_a, c51_d, c50_r, c50_a, c50_d);
  BrzSequence_2_s1_S I510 (c45_r, c45_a, c46_r, c46_a, c47_r, c47_a);
  BrzFetch_33_s5_false I511 (c46_r, c46_a, c43_r, c43_a, c43_d, c48_r, c48_a, c48_d);
  BrzFetch_33_s5_false I512 (c47_r, c47_a, c49_r, c49_a, c49_d, c44_r, c44_a, c44_d);
  BrzVariable_33_1_s0_ I513 (c48_r, c48_a, c48_d, c49_r, c49_a, c49_d);
  BrzCombine_33_32_1 I514 (c43_r, c43_a, c43_d, c42_r, c42_a, c42_d, c38_r, c38_a, c38_d);
  BrzSlice_32_34_1 I515 (c42_r, c42_a, c42_d, c41_r, c41_a, c41_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I516 (c41_r, c41_a, c41_d, c40_r, c40_a, c40_d, c39_r, c39_a, c39_d);
  BrzSlice_1_34_32 I517 (c38_r, c38_a, c38_d, c37_r, c37_a, c37_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I518 (c37_r, c37_a, c37_d, c36_r, c36_a, c36_d, c35_r, c35_a, c35_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I519 (c34_r, c34_a, c34_d, c33_r, c33_a, c33_d, c31_r, c31_a, c31_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I520 (c33_r, c33_a, c33_d, c32_r, c32_a, c32_d);
  BrzSequence_2_s1_S I521 (c26_r, c26_a, c27_r, c27_a, c28_r, c28_a);
  BrzFetch_33_s5_false I522 (c27_r, c27_a, c24_r, c24_a, c24_d, c29_r, c29_a, c29_d);
  BrzFetch_33_s5_false I523 (c28_r, c28_a, c30_r, c30_a, c30_d, c25_r, c25_a, c25_d);
  BrzVariable_33_1_s0_ I524 (c29_r, c29_a, c29_d, c30_r, c30_a, c30_d);
  BrzCombine_33_32_1 I525 (c24_r, c24_a, c24_d, c23_r, c23_a, c23_d, c19_r, c19_a, c19_d);
  BrzSlice_32_34_1 I526 (c23_r, c23_a, c23_d, c22_r, c22_a, c22_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I527 (c22_r, c22_a, c22_d, c21_r, c21_a, c21_d, c20_r, c20_a, c20_d);
  BrzSlice_1_34_32 I528 (c19_r, c19_a, c19_d, c18_r, c18_a, c18_d);
  BrzBinaryFunc_34_33_33_s3_Add_s4_true_s4_t_m2m I529 (c18_r, c18_a, c18_d, c17_r, c17_a, c17_d, c16_r, c16_a, c16_d);
  BrzSequence_2_s1_S I530 (c11_r, c11_a, c12_r, c12_a, c13_r, c13_a);
  BrzFetch_33_s5_false I531 (c12_r, c12_a, c9_r, c9_a, c9_d, c14_r, c14_a, c14_d);
  BrzFetch_33_s5_false I532 (c13_r, c13_a, c15_r, c15_a, c15_d, c10_r, c10_a, c10_d);
  BrzVariable_33_1_s0_ I533 (c14_r, c14_a, c14_d, c15_r, c15_a, c15_d);
  BrzCombine_33_32_1 I534 (c9_r, c9_a, c9_d, c8_r, c8_a, c8_d, c7_r, c7_a, c7_d);
  BrzFetch_32_s5_false I535 (c6_r, c6_a, c5_r, c5_a, c5_d, z_0r, z_0a, z_0d);
endmodule


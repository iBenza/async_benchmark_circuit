/*
    `booth_mul8.v'
    Balsa Verilog netlist file
    Created: Tue Jan 14 14:23:13 JST 2014
    By: xaos@kikurage (Linux)
    With net-verilog (balsa-netlist) version: 4.0
    Using technology: aclass/four_b_rb
    Command line : (balsa-netlist -Xaclass booth_mul8)

    Using `propagate-globals'
    The design contains no global nets
*/

module buf1 (
  z,
  a
);
  output z;
  input a;
  wire na_0n;
  IV I0 (z, na_0n);
  IV I1 (na_0n, a);
endmodule

module BrzAdapt_17_9_s5_false_s5_false (
  out_0r, out_0a, out_0d,
  inp_0r, inp_0a, inp_0d
);
  input out_0r;
  output out_0a;
  output [16:0] out_0d;
  output inp_0r;
  input inp_0a;
  input [8:0] inp_0d;
  wire extend_0n;
  wire gnd;
  GND gnd_cell_instance (gnd);
  assign out_0a = inp_0a;
  assign inp_0r = out_0r;
  assign out_0d[9] = gnd;
  assign out_0d[10] = gnd;
  assign out_0d[11] = gnd;
  assign out_0d[12] = gnd;
  assign out_0d[13] = gnd;
  assign out_0d[14] = gnd;
  assign out_0d[15] = gnd;
  assign out_0d[16] = gnd;
  assign out_0d[0] = inp_0d[0];
  assign out_0d[1] = inp_0d[1];
  assign out_0d[2] = inp_0d[2];
  assign out_0d[3] = inp_0d[3];
  assign out_0d[4] = inp_0d[4];
  assign out_0d[5] = inp_0d[5];
  assign out_0d[6] = inp_0d[6];
  assign out_0d[7] = inp_0d[7];
  assign out_0d[8] = inp_0d[8];
endmodule

module demux2 (
  i,
  o0,
  o1,
  s
);
  input i;
  output o0;
  output o1;
  input s;
  wire ns_0n;
  AN2 I0 (o1, i, s);
  AN2 I1 (o0, i, ns_0n);
  IV I2 (ns_0n, s);
endmodule

module BrzBar_2 (
  guard_0r, guard_0a, guard_0d,
  activate_0r, activate_0a,
  guardInput_0r, guardInput_0a, guardInput_0d,
  guardInput_1r, guardInput_1a, guardInput_1d,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a
);
  input guard_0r;
  output guard_0a;
  output guard_0d;
  input activate_0r;
  output activate_0a;
  output guardInput_0r;
  input guardInput_0a;
  input guardInput_0d;
  output guardInput_1r;
  input guardInput_1a;
  input guardInput_1d;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  wire [2:0] bypass_0n;
  wire [1:0] outReq_0n;
  C2 I0 (activateOut_0r, activate_0r, outReq_0n[0]);
  C2 I1 (activateOut_1r, activate_0r, outReq_0n[1]);
  demux2 I2 (bypass_0n[0], bypass_0n[1], outReq_0n[0], guardInput_0d);
  demux2 I3 (bypass_0n[1], bypass_0n[2], outReq_0n[1], guardInput_1d);
  assign bypass_0n[0] = activate_0r;
  OR3 I5 (activate_0a, activateOut_0a, activateOut_1a, bypass_0n[2]);
  OR2 I6 (guard_0d, guardInput_0d, guardInput_1d);
  C2 I7 (guard_0a, guardInput_0a, guardInput_1a);
  assign guardInput_0r = guard_0r;
  assign guardInput_1r = guard_0r;
endmodule

module BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m (
  out_0r, out_0a, out_0d,
  inpA_0r, inpA_0a, inpA_0d,
  inpB_0r, inpB_0a, inpB_0d
);
  input out_0r;
  output out_0a;
  output out_0d;
  output inpA_0r;
  input inpA_0a;
  input inpA_0d;
  output inpB_0r;
  input inpB_0a;
  input inpB_0d;
  wire start_0n;
  wire nStart_0n;
  wire [1:0] nCv_0n;
  wire [1:0] c_0n;
  wire eq_0n;
  wire addOut_0n;
  wire w_0n;
  wire n_0n;
  wire v_0n;
  wire z_0n;
  wire nz_0n;
  wire nxv_0n;
  wire done_0n;
  AN2 I0 (out_0d, n_0n, w_0n);
  assign done_0n = start_0n;
  assign n_0n = inpB_0d;
  assign w_0n = inpA_0d;
  assign out_0a = done_0n;
  C2 I5 (start_0n, inpA_0a, inpB_0a);
  assign inpA_0r = out_0r;
  assign inpB_0r = out_0r;
endmodule

module ao22 (
  q,
  i0,
  i1,
  i2,
  i3
);
  output q;
  input i0;
  input i1;
  input i2;
  input i3;
  wire [1:0] int_0n;
  OR2 I0 (q, int_0n[0], int_0n[1]);
  AN2 I1 (int_0n[1], i2, i3);
  AN2 I2 (int_0n[0], i0, i1);
endmodule

module mux2 (
  out,
  in0,
  in1,
  sel
);
  output out;
  input in0;
  input in1;
  input sel;
  wire nsel_0n;
  ao22 I0 (out, in0, nsel_0n, in1, sel);
  IV I1 (nsel_0n, sel);
endmodule

module aoi22 (
  q,
  i0,
  i1,
  i2,
  i3
);
  output q;
  input i0;
  input i1;
  input i2;
  input i3;
  wire [1:0] int_0n;
  NR2 I0 (q, int_0n[0], int_0n[1]);
  AN2 I1 (int_0n[1], i2, i3);
  AN2 I2 (int_0n[0], i0, i1);
endmodule

module nmux2 (
  out,
  in0,
  in1,
  sel
);
  output out;
  input in0;
  input in1;
  input sel;
  wire nsel_0n;
  aoi22 I0 (out, in0, nsel_0n, in1, sel);
  IV I1 (nsel_0n, sel);
endmodule

module balsa_fa (
  nStart,
  A,
  B,
  nCVi,
  Ci,
  nCVo,
  Co,
  sum
);
  input nStart;
  input A;
  input B;
  input nCVi;
  input Ci;
  output nCVo;
  output Co;
  output sum;
  wire start;
  wire ha;
  wire cv;
  IV I0 (start, nStart);
  NR2 I1 (cv, nStart, nCVi);
  nmux2 I2 (nCVo, start, cv, ha);
  mux2 I3 (Co, A, Ci, ha);
  EO I4 (ha, A, B);
  EO I5 (sum, ha, Ci);
endmodule

module BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m (
  out_0r, out_0a, out_0d,
  inpA_0r, inpA_0a, inpA_0d,
  inpB_0r, inpB_0a, inpB_0d
);
  input out_0r;
  output out_0a;
  output [17:0] out_0d;
  output inpA_0r;
  input inpA_0a;
  input [16:0] inpA_0d;
  output inpB_0r;
  input inpB_0a;
  input [16:0] inpB_0d;
  wire [6:0] internal_0n;
  wire start_0n;
  wire nStart_0n;
  wire [17:0] nCv_0n;
  wire [17:0] c_0n;
  wire [16:0] eq_0n;
  wire [16:0] addOut_0n;
  wire [16:0] w_0n;
  wire [16:0] n_0n;
  wire v_0n;
  wire z_0n;
  wire nz_0n;
  wire nxv_0n;
  wire done_0n;
  wire gnd;
  GND gnd_cell_instance (gnd);
  NR4 I0 (internal_0n[0], nCv_0n[1], nCv_0n[2], nCv_0n[3], nCv_0n[4]);
  NR4 I1 (internal_0n[1], nCv_0n[5], nCv_0n[6], nCv_0n[7], nCv_0n[8]);
  NR4 I2 (internal_0n[2], nCv_0n[9], nCv_0n[10], nCv_0n[11], nCv_0n[12]);
  NR2 I3 (internal_0n[3], nCv_0n[13], nCv_0n[14]);
  NR3 I4 (internal_0n[4], nCv_0n[15], nCv_0n[16], nCv_0n[17]);
  ND2 I5 (internal_0n[5], internal_0n[0], internal_0n[1]);
  ND3 I6 (internal_0n[6], internal_0n[2], internal_0n[3], internal_0n[4]);
  NR2 I7 (done_0n, internal_0n[5], internal_0n[6]);
  assign out_0d[0] = addOut_0n[0];
  assign out_0d[1] = addOut_0n[1];
  assign out_0d[2] = addOut_0n[2];
  assign out_0d[3] = addOut_0n[3];
  assign out_0d[4] = addOut_0n[4];
  assign out_0d[5] = addOut_0n[5];
  assign out_0d[6] = addOut_0n[6];
  assign out_0d[7] = addOut_0n[7];
  assign out_0d[8] = addOut_0n[8];
  assign out_0d[9] = addOut_0n[9];
  assign out_0d[10] = addOut_0n[10];
  assign out_0d[11] = addOut_0n[11];
  assign out_0d[12] = addOut_0n[12];
  assign out_0d[13] = addOut_0n[13];
  assign out_0d[14] = addOut_0n[14];
  assign out_0d[15] = addOut_0n[15];
  assign out_0d[16] = addOut_0n[16];
  assign out_0d[17] = c_0n[17];
  balsa_fa I26 (nStart_0n, n_0n[0], w_0n[0], nCv_0n[0], c_0n[0], nCv_0n[1], c_0n[1], addOut_0n[0]);
  balsa_fa I27 (nStart_0n, n_0n[1], w_0n[1], nCv_0n[1], c_0n[1], nCv_0n[2], c_0n[2], addOut_0n[1]);
  balsa_fa I28 (nStart_0n, n_0n[2], w_0n[2], nCv_0n[2], c_0n[2], nCv_0n[3], c_0n[3], addOut_0n[2]);
  balsa_fa I29 (nStart_0n, n_0n[3], w_0n[3], nCv_0n[3], c_0n[3], nCv_0n[4], c_0n[4], addOut_0n[3]);
  balsa_fa I30 (nStart_0n, n_0n[4], w_0n[4], nCv_0n[4], c_0n[4], nCv_0n[5], c_0n[5], addOut_0n[4]);
  balsa_fa I31 (nStart_0n, n_0n[5], w_0n[5], nCv_0n[5], c_0n[5], nCv_0n[6], c_0n[6], addOut_0n[5]);
  balsa_fa I32 (nStart_0n, n_0n[6], w_0n[6], nCv_0n[6], c_0n[6], nCv_0n[7], c_0n[7], addOut_0n[6]);
  balsa_fa I33 (nStart_0n, n_0n[7], w_0n[7], nCv_0n[7], c_0n[7], nCv_0n[8], c_0n[8], addOut_0n[7]);
  balsa_fa I34 (nStart_0n, n_0n[8], w_0n[8], nCv_0n[8], c_0n[8], nCv_0n[9], c_0n[9], addOut_0n[8]);
  balsa_fa I35 (nStart_0n, n_0n[9], w_0n[9], nCv_0n[9], c_0n[9], nCv_0n[10], c_0n[10], addOut_0n[9]);
  balsa_fa I36 (nStart_0n, n_0n[10], w_0n[10], nCv_0n[10], c_0n[10], nCv_0n[11], c_0n[11], addOut_0n[10]);
  balsa_fa I37 (nStart_0n, n_0n[11], w_0n[11], nCv_0n[11], c_0n[11], nCv_0n[12], c_0n[12], addOut_0n[11]);
  balsa_fa I38 (nStart_0n, n_0n[12], w_0n[12], nCv_0n[12], c_0n[12], nCv_0n[13], c_0n[13], addOut_0n[12]);
  balsa_fa I39 (nStart_0n, n_0n[13], w_0n[13], nCv_0n[13], c_0n[13], nCv_0n[14], c_0n[14], addOut_0n[13]);
  balsa_fa I40 (nStart_0n, n_0n[14], w_0n[14], nCv_0n[14], c_0n[14], nCv_0n[15], c_0n[15], addOut_0n[14]);
  balsa_fa I41 (nStart_0n, n_0n[15], w_0n[15], nCv_0n[15], c_0n[15], nCv_0n[16], c_0n[16], addOut_0n[15]);
  balsa_fa I42 (nStart_0n, n_0n[16], w_0n[16], nCv_0n[16], c_0n[16], nCv_0n[17], c_0n[17], addOut_0n[16]);
  assign nCv_0n[0] = nStart_0n;
  assign c_0n[0] = gnd;
  IV I45 (nStart_0n, start_0n);
  assign n_0n[0] = inpB_0d[0];
  assign n_0n[1] = inpB_0d[1];
  assign n_0n[2] = inpB_0d[2];
  assign n_0n[3] = inpB_0d[3];
  assign n_0n[4] = inpB_0d[4];
  assign n_0n[5] = inpB_0d[5];
  assign n_0n[6] = inpB_0d[6];
  assign n_0n[7] = inpB_0d[7];
  assign n_0n[8] = inpB_0d[8];
  assign n_0n[9] = inpB_0d[9];
  assign n_0n[10] = inpB_0d[10];
  assign n_0n[11] = inpB_0d[11];
  assign n_0n[12] = inpB_0d[12];
  assign n_0n[13] = inpB_0d[13];
  assign n_0n[14] = inpB_0d[14];
  assign n_0n[15] = inpB_0d[15];
  assign n_0n[16] = inpB_0d[16];
  assign w_0n[0] = inpA_0d[0];
  assign w_0n[1] = inpA_0d[1];
  assign w_0n[2] = inpA_0d[2];
  assign w_0n[3] = inpA_0d[3];
  assign w_0n[4] = inpA_0d[4];
  assign w_0n[5] = inpA_0d[5];
  assign w_0n[6] = inpA_0d[6];
  assign w_0n[7] = inpA_0d[7];
  assign w_0n[8] = inpA_0d[8];
  assign w_0n[9] = inpA_0d[9];
  assign w_0n[10] = inpA_0d[10];
  assign w_0n[11] = inpA_0d[11];
  assign w_0n[12] = inpA_0d[12];
  assign w_0n[13] = inpA_0d[13];
  assign w_0n[14] = inpA_0d[14];
  assign w_0n[15] = inpA_0d[15];
  assign w_0n[16] = inpA_0d[16];
  assign out_0a = done_0n;
  C2 I81 (start_0n, inpA_0a, inpB_0a);
  assign inpA_0r = out_0r;
  assign inpB_0r = out_0r;
endmodule

module BrzCallMux_17_25 (
  inp_0r, inp_0a, inp_0d,
  inp_1r, inp_1a, inp_1d,
  inp_2r, inp_2a, inp_2d,
  inp_3r, inp_3a, inp_3d,
  inp_4r, inp_4a, inp_4d,
  inp_5r, inp_5a, inp_5d,
  inp_6r, inp_6a, inp_6d,
  inp_7r, inp_7a, inp_7d,
  inp_8r, inp_8a, inp_8d,
  inp_9r, inp_9a, inp_9d,
  inp_10r, inp_10a, inp_10d,
  inp_11r, inp_11a, inp_11d,
  inp_12r, inp_12a, inp_12d,
  inp_13r, inp_13a, inp_13d,
  inp_14r, inp_14a, inp_14d,
  inp_15r, inp_15a, inp_15d,
  inp_16r, inp_16a, inp_16d,
  inp_17r, inp_17a, inp_17d,
  inp_18r, inp_18a, inp_18d,
  inp_19r, inp_19a, inp_19d,
  inp_20r, inp_20a, inp_20d,
  inp_21r, inp_21a, inp_21d,
  inp_22r, inp_22a, inp_22d,
  inp_23r, inp_23a, inp_23d,
  inp_24r, inp_24a, inp_24d,
  out_0r, out_0a, out_0d
);
  input inp_0r;
  output inp_0a;
  input [16:0] inp_0d;
  input inp_1r;
  output inp_1a;
  input [16:0] inp_1d;
  input inp_2r;
  output inp_2a;
  input [16:0] inp_2d;
  input inp_3r;
  output inp_3a;
  input [16:0] inp_3d;
  input inp_4r;
  output inp_4a;
  input [16:0] inp_4d;
  input inp_5r;
  output inp_5a;
  input [16:0] inp_5d;
  input inp_6r;
  output inp_6a;
  input [16:0] inp_6d;
  input inp_7r;
  output inp_7a;
  input [16:0] inp_7d;
  input inp_8r;
  output inp_8a;
  input [16:0] inp_8d;
  input inp_9r;
  output inp_9a;
  input [16:0] inp_9d;
  input inp_10r;
  output inp_10a;
  input [16:0] inp_10d;
  input inp_11r;
  output inp_11a;
  input [16:0] inp_11d;
  input inp_12r;
  output inp_12a;
  input [16:0] inp_12d;
  input inp_13r;
  output inp_13a;
  input [16:0] inp_13d;
  input inp_14r;
  output inp_14a;
  input [16:0] inp_14d;
  input inp_15r;
  output inp_15a;
  input [16:0] inp_15d;
  input inp_16r;
  output inp_16a;
  input [16:0] inp_16d;
  input inp_17r;
  output inp_17a;
  input [16:0] inp_17d;
  input inp_18r;
  output inp_18a;
  input [16:0] inp_18d;
  input inp_19r;
  output inp_19a;
  input [16:0] inp_19d;
  input inp_20r;
  output inp_20a;
  input [16:0] inp_20d;
  input inp_21r;
  output inp_21a;
  input [16:0] inp_21d;
  input inp_22r;
  output inp_22a;
  input [16:0] inp_22d;
  input inp_23r;
  output inp_23a;
  input [16:0] inp_23d;
  input inp_24r;
  output inp_24a;
  input [16:0] inp_24d;
  output out_0r;
  input out_0a;
  output [16:0] out_0d;
  wire [161:0] internal_0n;
  wire [16:0] muxOut_0n;
  wire select_0n;
  wire nselect_0n;
  wire [24:0] nwaySelect_0n;
  wire [16:0] nwayMuxOut_0n;
  wire [16:0] nwayMuxOut_1n;
  wire [16:0] nwayMuxOut_2n;
  wire [16:0] nwayMuxOut_3n;
  wire [16:0] nwayMuxOut_4n;
  wire [16:0] nwayMuxOut_5n;
  wire [16:0] nwayMuxOut_6n;
  wire [16:0] nwayMuxOut_7n;
  wire [16:0] nwayMuxOut_8n;
  wire [16:0] nwayMuxOut_9n;
  wire [16:0] nwayMuxOut_10n;
  wire [16:0] nwayMuxOut_11n;
  wire [16:0] nwayMuxOut_12n;
  wire [16:0] nwayMuxOut_13n;
  wire [16:0] nwayMuxOut_14n;
  wire [16:0] nwayMuxOut_15n;
  wire [16:0] nwayMuxOut_16n;
  wire [16:0] nwayMuxOut_17n;
  wire [16:0] nwayMuxOut_18n;
  wire [16:0] nwayMuxOut_19n;
  wire [16:0] nwayMuxOut_20n;
  wire [16:0] nwayMuxOut_21n;
  wire [16:0] nwayMuxOut_22n;
  wire [16:0] nwayMuxOut_23n;
  wire [16:0] nwayMuxOut_24n;
  ND4 I0 (internal_0n[0], nwayMuxOut_0n[0], nwayMuxOut_1n[0], nwayMuxOut_2n[0], nwayMuxOut_3n[0]);
  ND4 I1 (internal_0n[1], nwayMuxOut_4n[0], nwayMuxOut_5n[0], nwayMuxOut_6n[0], nwayMuxOut_7n[0]);
  ND4 I2 (internal_0n[2], nwayMuxOut_8n[0], nwayMuxOut_9n[0], nwayMuxOut_10n[0], nwayMuxOut_11n[0]);
  ND4 I3 (internal_0n[3], nwayMuxOut_12n[0], nwayMuxOut_13n[0], nwayMuxOut_14n[0], nwayMuxOut_15n[0]);
  ND4 I4 (internal_0n[4], nwayMuxOut_16n[0], nwayMuxOut_17n[0], nwayMuxOut_18n[0], nwayMuxOut_19n[0]);
  ND2 I5 (internal_0n[5], nwayMuxOut_20n[0], nwayMuxOut_21n[0]);
  ND3 I6 (internal_0n[6], nwayMuxOut_22n[0], nwayMuxOut_23n[0], nwayMuxOut_24n[0]);
  NR4 I7 (internal_0n[7], internal_0n[0], internal_0n[1], internal_0n[2], internal_0n[3]);
  NR3 I8 (internal_0n[8], internal_0n[4], internal_0n[5], internal_0n[6]);
  ND2 I9 (out_0d[0], internal_0n[7], internal_0n[8]);
  ND4 I10 (internal_0n[9], nwayMuxOut_0n[1], nwayMuxOut_1n[1], nwayMuxOut_2n[1], nwayMuxOut_3n[1]);
  ND4 I11 (internal_0n[10], nwayMuxOut_4n[1], nwayMuxOut_5n[1], nwayMuxOut_6n[1], nwayMuxOut_7n[1]);
  ND4 I12 (internal_0n[11], nwayMuxOut_8n[1], nwayMuxOut_9n[1], nwayMuxOut_10n[1], nwayMuxOut_11n[1]);
  ND4 I13 (internal_0n[12], nwayMuxOut_12n[1], nwayMuxOut_13n[1], nwayMuxOut_14n[1], nwayMuxOut_15n[1]);
  ND4 I14 (internal_0n[13], nwayMuxOut_16n[1], nwayMuxOut_17n[1], nwayMuxOut_18n[1], nwayMuxOut_19n[1]);
  ND2 I15 (internal_0n[14], nwayMuxOut_20n[1], nwayMuxOut_21n[1]);
  ND3 I16 (internal_0n[15], nwayMuxOut_22n[1], nwayMuxOut_23n[1], nwayMuxOut_24n[1]);
  NR4 I17 (internal_0n[16], internal_0n[9], internal_0n[10], internal_0n[11], internal_0n[12]);
  NR3 I18 (internal_0n[17], internal_0n[13], internal_0n[14], internal_0n[15]);
  ND2 I19 (out_0d[1], internal_0n[16], internal_0n[17]);
  ND4 I20 (internal_0n[18], nwayMuxOut_0n[2], nwayMuxOut_1n[2], nwayMuxOut_2n[2], nwayMuxOut_3n[2]);
  ND4 I21 (internal_0n[19], nwayMuxOut_4n[2], nwayMuxOut_5n[2], nwayMuxOut_6n[2], nwayMuxOut_7n[2]);
  ND4 I22 (internal_0n[20], nwayMuxOut_8n[2], nwayMuxOut_9n[2], nwayMuxOut_10n[2], nwayMuxOut_11n[2]);
  ND4 I23 (internal_0n[21], nwayMuxOut_12n[2], nwayMuxOut_13n[2], nwayMuxOut_14n[2], nwayMuxOut_15n[2]);
  ND4 I24 (internal_0n[22], nwayMuxOut_16n[2], nwayMuxOut_17n[2], nwayMuxOut_18n[2], nwayMuxOut_19n[2]);
  ND2 I25 (internal_0n[23], nwayMuxOut_20n[2], nwayMuxOut_21n[2]);
  ND3 I26 (internal_0n[24], nwayMuxOut_22n[2], nwayMuxOut_23n[2], nwayMuxOut_24n[2]);
  NR4 I27 (internal_0n[25], internal_0n[18], internal_0n[19], internal_0n[20], internal_0n[21]);
  NR3 I28 (internal_0n[26], internal_0n[22], internal_0n[23], internal_0n[24]);
  ND2 I29 (out_0d[2], internal_0n[25], internal_0n[26]);
  ND4 I30 (internal_0n[27], nwayMuxOut_0n[3], nwayMuxOut_1n[3], nwayMuxOut_2n[3], nwayMuxOut_3n[3]);
  ND4 I31 (internal_0n[28], nwayMuxOut_4n[3], nwayMuxOut_5n[3], nwayMuxOut_6n[3], nwayMuxOut_7n[3]);
  ND4 I32 (internal_0n[29], nwayMuxOut_8n[3], nwayMuxOut_9n[3], nwayMuxOut_10n[3], nwayMuxOut_11n[3]);
  ND4 I33 (internal_0n[30], nwayMuxOut_12n[3], nwayMuxOut_13n[3], nwayMuxOut_14n[3], nwayMuxOut_15n[3]);
  ND4 I34 (internal_0n[31], nwayMuxOut_16n[3], nwayMuxOut_17n[3], nwayMuxOut_18n[3], nwayMuxOut_19n[3]);
  ND2 I35 (internal_0n[32], nwayMuxOut_20n[3], nwayMuxOut_21n[3]);
  ND3 I36 (internal_0n[33], nwayMuxOut_22n[3], nwayMuxOut_23n[3], nwayMuxOut_24n[3]);
  NR4 I37 (internal_0n[34], internal_0n[27], internal_0n[28], internal_0n[29], internal_0n[30]);
  NR3 I38 (internal_0n[35], internal_0n[31], internal_0n[32], internal_0n[33]);
  ND2 I39 (out_0d[3], internal_0n[34], internal_0n[35]);
  ND4 I40 (internal_0n[36], nwayMuxOut_0n[4], nwayMuxOut_1n[4], nwayMuxOut_2n[4], nwayMuxOut_3n[4]);
  ND4 I41 (internal_0n[37], nwayMuxOut_4n[4], nwayMuxOut_5n[4], nwayMuxOut_6n[4], nwayMuxOut_7n[4]);
  ND4 I42 (internal_0n[38], nwayMuxOut_8n[4], nwayMuxOut_9n[4], nwayMuxOut_10n[4], nwayMuxOut_11n[4]);
  ND4 I43 (internal_0n[39], nwayMuxOut_12n[4], nwayMuxOut_13n[4], nwayMuxOut_14n[4], nwayMuxOut_15n[4]);
  ND4 I44 (internal_0n[40], nwayMuxOut_16n[4], nwayMuxOut_17n[4], nwayMuxOut_18n[4], nwayMuxOut_19n[4]);
  ND2 I45 (internal_0n[41], nwayMuxOut_20n[4], nwayMuxOut_21n[4]);
  ND3 I46 (internal_0n[42], nwayMuxOut_22n[4], nwayMuxOut_23n[4], nwayMuxOut_24n[4]);
  NR4 I47 (internal_0n[43], internal_0n[36], internal_0n[37], internal_0n[38], internal_0n[39]);
  NR3 I48 (internal_0n[44], internal_0n[40], internal_0n[41], internal_0n[42]);
  ND2 I49 (out_0d[4], internal_0n[43], internal_0n[44]);
  ND4 I50 (internal_0n[45], nwayMuxOut_0n[5], nwayMuxOut_1n[5], nwayMuxOut_2n[5], nwayMuxOut_3n[5]);
  ND4 I51 (internal_0n[46], nwayMuxOut_4n[5], nwayMuxOut_5n[5], nwayMuxOut_6n[5], nwayMuxOut_7n[5]);
  ND4 I52 (internal_0n[47], nwayMuxOut_8n[5], nwayMuxOut_9n[5], nwayMuxOut_10n[5], nwayMuxOut_11n[5]);
  ND4 I53 (internal_0n[48], nwayMuxOut_12n[5], nwayMuxOut_13n[5], nwayMuxOut_14n[5], nwayMuxOut_15n[5]);
  ND4 I54 (internal_0n[49], nwayMuxOut_16n[5], nwayMuxOut_17n[5], nwayMuxOut_18n[5], nwayMuxOut_19n[5]);
  ND2 I55 (internal_0n[50], nwayMuxOut_20n[5], nwayMuxOut_21n[5]);
  ND3 I56 (internal_0n[51], nwayMuxOut_22n[5], nwayMuxOut_23n[5], nwayMuxOut_24n[5]);
  NR4 I57 (internal_0n[52], internal_0n[45], internal_0n[46], internal_0n[47], internal_0n[48]);
  NR3 I58 (internal_0n[53], internal_0n[49], internal_0n[50], internal_0n[51]);
  ND2 I59 (out_0d[5], internal_0n[52], internal_0n[53]);
  ND4 I60 (internal_0n[54], nwayMuxOut_0n[6], nwayMuxOut_1n[6], nwayMuxOut_2n[6], nwayMuxOut_3n[6]);
  ND4 I61 (internal_0n[55], nwayMuxOut_4n[6], nwayMuxOut_5n[6], nwayMuxOut_6n[6], nwayMuxOut_7n[6]);
  ND4 I62 (internal_0n[56], nwayMuxOut_8n[6], nwayMuxOut_9n[6], nwayMuxOut_10n[6], nwayMuxOut_11n[6]);
  ND4 I63 (internal_0n[57], nwayMuxOut_12n[6], nwayMuxOut_13n[6], nwayMuxOut_14n[6], nwayMuxOut_15n[6]);
  ND4 I64 (internal_0n[58], nwayMuxOut_16n[6], nwayMuxOut_17n[6], nwayMuxOut_18n[6], nwayMuxOut_19n[6]);
  ND2 I65 (internal_0n[59], nwayMuxOut_20n[6], nwayMuxOut_21n[6]);
  ND3 I66 (internal_0n[60], nwayMuxOut_22n[6], nwayMuxOut_23n[6], nwayMuxOut_24n[6]);
  NR4 I67 (internal_0n[61], internal_0n[54], internal_0n[55], internal_0n[56], internal_0n[57]);
  NR3 I68 (internal_0n[62], internal_0n[58], internal_0n[59], internal_0n[60]);
  ND2 I69 (out_0d[6], internal_0n[61], internal_0n[62]);
  ND4 I70 (internal_0n[63], nwayMuxOut_0n[7], nwayMuxOut_1n[7], nwayMuxOut_2n[7], nwayMuxOut_3n[7]);
  ND4 I71 (internal_0n[64], nwayMuxOut_4n[7], nwayMuxOut_5n[7], nwayMuxOut_6n[7], nwayMuxOut_7n[7]);
  ND4 I72 (internal_0n[65], nwayMuxOut_8n[7], nwayMuxOut_9n[7], nwayMuxOut_10n[7], nwayMuxOut_11n[7]);
  ND4 I73 (internal_0n[66], nwayMuxOut_12n[7], nwayMuxOut_13n[7], nwayMuxOut_14n[7], nwayMuxOut_15n[7]);
  ND4 I74 (internal_0n[67], nwayMuxOut_16n[7], nwayMuxOut_17n[7], nwayMuxOut_18n[7], nwayMuxOut_19n[7]);
  ND2 I75 (internal_0n[68], nwayMuxOut_20n[7], nwayMuxOut_21n[7]);
  ND3 I76 (internal_0n[69], nwayMuxOut_22n[7], nwayMuxOut_23n[7], nwayMuxOut_24n[7]);
  NR4 I77 (internal_0n[70], internal_0n[63], internal_0n[64], internal_0n[65], internal_0n[66]);
  NR3 I78 (internal_0n[71], internal_0n[67], internal_0n[68], internal_0n[69]);
  ND2 I79 (out_0d[7], internal_0n[70], internal_0n[71]);
  ND4 I80 (internal_0n[72], nwayMuxOut_0n[8], nwayMuxOut_1n[8], nwayMuxOut_2n[8], nwayMuxOut_3n[8]);
  ND4 I81 (internal_0n[73], nwayMuxOut_4n[8], nwayMuxOut_5n[8], nwayMuxOut_6n[8], nwayMuxOut_7n[8]);
  ND4 I82 (internal_0n[74], nwayMuxOut_8n[8], nwayMuxOut_9n[8], nwayMuxOut_10n[8], nwayMuxOut_11n[8]);
  ND4 I83 (internal_0n[75], nwayMuxOut_12n[8], nwayMuxOut_13n[8], nwayMuxOut_14n[8], nwayMuxOut_15n[8]);
  ND4 I84 (internal_0n[76], nwayMuxOut_16n[8], nwayMuxOut_17n[8], nwayMuxOut_18n[8], nwayMuxOut_19n[8]);
  ND2 I85 (internal_0n[77], nwayMuxOut_20n[8], nwayMuxOut_21n[8]);
  ND3 I86 (internal_0n[78], nwayMuxOut_22n[8], nwayMuxOut_23n[8], nwayMuxOut_24n[8]);
  NR4 I87 (internal_0n[79], internal_0n[72], internal_0n[73], internal_0n[74], internal_0n[75]);
  NR3 I88 (internal_0n[80], internal_0n[76], internal_0n[77], internal_0n[78]);
  ND2 I89 (out_0d[8], internal_0n[79], internal_0n[80]);
  ND4 I90 (internal_0n[81], nwayMuxOut_0n[9], nwayMuxOut_1n[9], nwayMuxOut_2n[9], nwayMuxOut_3n[9]);
  ND4 I91 (internal_0n[82], nwayMuxOut_4n[9], nwayMuxOut_5n[9], nwayMuxOut_6n[9], nwayMuxOut_7n[9]);
  ND4 I92 (internal_0n[83], nwayMuxOut_8n[9], nwayMuxOut_9n[9], nwayMuxOut_10n[9], nwayMuxOut_11n[9]);
  ND4 I93 (internal_0n[84], nwayMuxOut_12n[9], nwayMuxOut_13n[9], nwayMuxOut_14n[9], nwayMuxOut_15n[9]);
  ND4 I94 (internal_0n[85], nwayMuxOut_16n[9], nwayMuxOut_17n[9], nwayMuxOut_18n[9], nwayMuxOut_19n[9]);
  ND2 I95 (internal_0n[86], nwayMuxOut_20n[9], nwayMuxOut_21n[9]);
  ND3 I96 (internal_0n[87], nwayMuxOut_22n[9], nwayMuxOut_23n[9], nwayMuxOut_24n[9]);
  NR4 I97 (internal_0n[88], internal_0n[81], internal_0n[82], internal_0n[83], internal_0n[84]);
  NR3 I98 (internal_0n[89], internal_0n[85], internal_0n[86], internal_0n[87]);
  ND2 I99 (out_0d[9], internal_0n[88], internal_0n[89]);
  ND4 I100 (internal_0n[90], nwayMuxOut_0n[10], nwayMuxOut_1n[10], nwayMuxOut_2n[10], nwayMuxOut_3n[10]);
  ND4 I101 (internal_0n[91], nwayMuxOut_4n[10], nwayMuxOut_5n[10], nwayMuxOut_6n[10], nwayMuxOut_7n[10]);
  ND4 I102 (internal_0n[92], nwayMuxOut_8n[10], nwayMuxOut_9n[10], nwayMuxOut_10n[10], nwayMuxOut_11n[10]);
  ND4 I103 (internal_0n[93], nwayMuxOut_12n[10], nwayMuxOut_13n[10], nwayMuxOut_14n[10], nwayMuxOut_15n[10]);
  ND4 I104 (internal_0n[94], nwayMuxOut_16n[10], nwayMuxOut_17n[10], nwayMuxOut_18n[10], nwayMuxOut_19n[10]);
  ND2 I105 (internal_0n[95], nwayMuxOut_20n[10], nwayMuxOut_21n[10]);
  ND3 I106 (internal_0n[96], nwayMuxOut_22n[10], nwayMuxOut_23n[10], nwayMuxOut_24n[10]);
  NR4 I107 (internal_0n[97], internal_0n[90], internal_0n[91], internal_0n[92], internal_0n[93]);
  NR3 I108 (internal_0n[98], internal_0n[94], internal_0n[95], internal_0n[96]);
  ND2 I109 (out_0d[10], internal_0n[97], internal_0n[98]);
  ND4 I110 (internal_0n[99], nwayMuxOut_0n[11], nwayMuxOut_1n[11], nwayMuxOut_2n[11], nwayMuxOut_3n[11]);
  ND4 I111 (internal_0n[100], nwayMuxOut_4n[11], nwayMuxOut_5n[11], nwayMuxOut_6n[11], nwayMuxOut_7n[11]);
  ND4 I112 (internal_0n[101], nwayMuxOut_8n[11], nwayMuxOut_9n[11], nwayMuxOut_10n[11], nwayMuxOut_11n[11]);
  ND4 I113 (internal_0n[102], nwayMuxOut_12n[11], nwayMuxOut_13n[11], nwayMuxOut_14n[11], nwayMuxOut_15n[11]);
  ND4 I114 (internal_0n[103], nwayMuxOut_16n[11], nwayMuxOut_17n[11], nwayMuxOut_18n[11], nwayMuxOut_19n[11]);
  ND2 I115 (internal_0n[104], nwayMuxOut_20n[11], nwayMuxOut_21n[11]);
  ND3 I116 (internal_0n[105], nwayMuxOut_22n[11], nwayMuxOut_23n[11], nwayMuxOut_24n[11]);
  NR4 I117 (internal_0n[106], internal_0n[99], internal_0n[100], internal_0n[101], internal_0n[102]);
  NR3 I118 (internal_0n[107], internal_0n[103], internal_0n[104], internal_0n[105]);
  ND2 I119 (out_0d[11], internal_0n[106], internal_0n[107]);
  ND4 I120 (internal_0n[108], nwayMuxOut_0n[12], nwayMuxOut_1n[12], nwayMuxOut_2n[12], nwayMuxOut_3n[12]);
  ND4 I121 (internal_0n[109], nwayMuxOut_4n[12], nwayMuxOut_5n[12], nwayMuxOut_6n[12], nwayMuxOut_7n[12]);
  ND4 I122 (internal_0n[110], nwayMuxOut_8n[12], nwayMuxOut_9n[12], nwayMuxOut_10n[12], nwayMuxOut_11n[12]);
  ND4 I123 (internal_0n[111], nwayMuxOut_12n[12], nwayMuxOut_13n[12], nwayMuxOut_14n[12], nwayMuxOut_15n[12]);
  ND4 I124 (internal_0n[112], nwayMuxOut_16n[12], nwayMuxOut_17n[12], nwayMuxOut_18n[12], nwayMuxOut_19n[12]);
  ND2 I125 (internal_0n[113], nwayMuxOut_20n[12], nwayMuxOut_21n[12]);
  ND3 I126 (internal_0n[114], nwayMuxOut_22n[12], nwayMuxOut_23n[12], nwayMuxOut_24n[12]);
  NR4 I127 (internal_0n[115], internal_0n[108], internal_0n[109], internal_0n[110], internal_0n[111]);
  NR3 I128 (internal_0n[116], internal_0n[112], internal_0n[113], internal_0n[114]);
  ND2 I129 (out_0d[12], internal_0n[115], internal_0n[116]);
  ND4 I130 (internal_0n[117], nwayMuxOut_0n[13], nwayMuxOut_1n[13], nwayMuxOut_2n[13], nwayMuxOut_3n[13]);
  ND4 I131 (internal_0n[118], nwayMuxOut_4n[13], nwayMuxOut_5n[13], nwayMuxOut_6n[13], nwayMuxOut_7n[13]);
  ND4 I132 (internal_0n[119], nwayMuxOut_8n[13], nwayMuxOut_9n[13], nwayMuxOut_10n[13], nwayMuxOut_11n[13]);
  ND4 I133 (internal_0n[120], nwayMuxOut_12n[13], nwayMuxOut_13n[13], nwayMuxOut_14n[13], nwayMuxOut_15n[13]);
  ND4 I134 (internal_0n[121], nwayMuxOut_16n[13], nwayMuxOut_17n[13], nwayMuxOut_18n[13], nwayMuxOut_19n[13]);
  ND2 I135 (internal_0n[122], nwayMuxOut_20n[13], nwayMuxOut_21n[13]);
  ND3 I136 (internal_0n[123], nwayMuxOut_22n[13], nwayMuxOut_23n[13], nwayMuxOut_24n[13]);
  NR4 I137 (internal_0n[124], internal_0n[117], internal_0n[118], internal_0n[119], internal_0n[120]);
  NR3 I138 (internal_0n[125], internal_0n[121], internal_0n[122], internal_0n[123]);
  ND2 I139 (out_0d[13], internal_0n[124], internal_0n[125]);
  ND4 I140 (internal_0n[126], nwayMuxOut_0n[14], nwayMuxOut_1n[14], nwayMuxOut_2n[14], nwayMuxOut_3n[14]);
  ND4 I141 (internal_0n[127], nwayMuxOut_4n[14], nwayMuxOut_5n[14], nwayMuxOut_6n[14], nwayMuxOut_7n[14]);
  ND4 I142 (internal_0n[128], nwayMuxOut_8n[14], nwayMuxOut_9n[14], nwayMuxOut_10n[14], nwayMuxOut_11n[14]);
  ND4 I143 (internal_0n[129], nwayMuxOut_12n[14], nwayMuxOut_13n[14], nwayMuxOut_14n[14], nwayMuxOut_15n[14]);
  ND4 I144 (internal_0n[130], nwayMuxOut_16n[14], nwayMuxOut_17n[14], nwayMuxOut_18n[14], nwayMuxOut_19n[14]);
  ND2 I145 (internal_0n[131], nwayMuxOut_20n[14], nwayMuxOut_21n[14]);
  ND3 I146 (internal_0n[132], nwayMuxOut_22n[14], nwayMuxOut_23n[14], nwayMuxOut_24n[14]);
  NR4 I147 (internal_0n[133], internal_0n[126], internal_0n[127], internal_0n[128], internal_0n[129]);
  NR3 I148 (internal_0n[134], internal_0n[130], internal_0n[131], internal_0n[132]);
  ND2 I149 (out_0d[14], internal_0n[133], internal_0n[134]);
  ND4 I150 (internal_0n[135], nwayMuxOut_0n[15], nwayMuxOut_1n[15], nwayMuxOut_2n[15], nwayMuxOut_3n[15]);
  ND4 I151 (internal_0n[136], nwayMuxOut_4n[15], nwayMuxOut_5n[15], nwayMuxOut_6n[15], nwayMuxOut_7n[15]);
  ND4 I152 (internal_0n[137], nwayMuxOut_8n[15], nwayMuxOut_9n[15], nwayMuxOut_10n[15], nwayMuxOut_11n[15]);
  ND4 I153 (internal_0n[138], nwayMuxOut_12n[15], nwayMuxOut_13n[15], nwayMuxOut_14n[15], nwayMuxOut_15n[15]);
  ND4 I154 (internal_0n[139], nwayMuxOut_16n[15], nwayMuxOut_17n[15], nwayMuxOut_18n[15], nwayMuxOut_19n[15]);
  ND2 I155 (internal_0n[140], nwayMuxOut_20n[15], nwayMuxOut_21n[15]);
  ND3 I156 (internal_0n[141], nwayMuxOut_22n[15], nwayMuxOut_23n[15], nwayMuxOut_24n[15]);
  NR4 I157 (internal_0n[142], internal_0n[135], internal_0n[136], internal_0n[137], internal_0n[138]);
  NR3 I158 (internal_0n[143], internal_0n[139], internal_0n[140], internal_0n[141]);
  ND2 I159 (out_0d[15], internal_0n[142], internal_0n[143]);
  ND4 I160 (internal_0n[144], nwayMuxOut_0n[16], nwayMuxOut_1n[16], nwayMuxOut_2n[16], nwayMuxOut_3n[16]);
  ND4 I161 (internal_0n[145], nwayMuxOut_4n[16], nwayMuxOut_5n[16], nwayMuxOut_6n[16], nwayMuxOut_7n[16]);
  ND4 I162 (internal_0n[146], nwayMuxOut_8n[16], nwayMuxOut_9n[16], nwayMuxOut_10n[16], nwayMuxOut_11n[16]);
  ND4 I163 (internal_0n[147], nwayMuxOut_12n[16], nwayMuxOut_13n[16], nwayMuxOut_14n[16], nwayMuxOut_15n[16]);
  ND4 I164 (internal_0n[148], nwayMuxOut_16n[16], nwayMuxOut_17n[16], nwayMuxOut_18n[16], nwayMuxOut_19n[16]);
  ND2 I165 (internal_0n[149], nwayMuxOut_20n[16], nwayMuxOut_21n[16]);
  ND3 I166 (internal_0n[150], nwayMuxOut_22n[16], nwayMuxOut_23n[16], nwayMuxOut_24n[16]);
  NR4 I167 (internal_0n[151], internal_0n[144], internal_0n[145], internal_0n[146], internal_0n[147]);
  NR3 I168 (internal_0n[152], internal_0n[148], internal_0n[149], internal_0n[150]);
  ND2 I169 (out_0d[16], internal_0n[151], internal_0n[152]);
  ND2 I170 (nwayMuxOut_0n[0], inp_0d[0], nwaySelect_0n[0]);
  ND2 I171 (nwayMuxOut_0n[1], inp_0d[1], nwaySelect_0n[0]);
  ND2 I172 (nwayMuxOut_0n[2], inp_0d[2], nwaySelect_0n[0]);
  ND2 I173 (nwayMuxOut_0n[3], inp_0d[3], nwaySelect_0n[0]);
  ND2 I174 (nwayMuxOut_0n[4], inp_0d[4], nwaySelect_0n[0]);
  ND2 I175 (nwayMuxOut_0n[5], inp_0d[5], nwaySelect_0n[0]);
  ND2 I176 (nwayMuxOut_0n[6], inp_0d[6], nwaySelect_0n[0]);
  ND2 I177 (nwayMuxOut_0n[7], inp_0d[7], nwaySelect_0n[0]);
  ND2 I178 (nwayMuxOut_0n[8], inp_0d[8], nwaySelect_0n[0]);
  ND2 I179 (nwayMuxOut_0n[9], inp_0d[9], nwaySelect_0n[0]);
  ND2 I180 (nwayMuxOut_0n[10], inp_0d[10], nwaySelect_0n[0]);
  ND2 I181 (nwayMuxOut_0n[11], inp_0d[11], nwaySelect_0n[0]);
  ND2 I182 (nwayMuxOut_0n[12], inp_0d[12], nwaySelect_0n[0]);
  ND2 I183 (nwayMuxOut_0n[13], inp_0d[13], nwaySelect_0n[0]);
  ND2 I184 (nwayMuxOut_0n[14], inp_0d[14], nwaySelect_0n[0]);
  ND2 I185 (nwayMuxOut_0n[15], inp_0d[15], nwaySelect_0n[0]);
  ND2 I186 (nwayMuxOut_0n[16], inp_0d[16], nwaySelect_0n[0]);
  ND2 I187 (nwayMuxOut_1n[0], inp_1d[0], nwaySelect_0n[1]);
  ND2 I188 (nwayMuxOut_1n[1], inp_1d[1], nwaySelect_0n[1]);
  ND2 I189 (nwayMuxOut_1n[2], inp_1d[2], nwaySelect_0n[1]);
  ND2 I190 (nwayMuxOut_1n[3], inp_1d[3], nwaySelect_0n[1]);
  ND2 I191 (nwayMuxOut_1n[4], inp_1d[4], nwaySelect_0n[1]);
  ND2 I192 (nwayMuxOut_1n[5], inp_1d[5], nwaySelect_0n[1]);
  ND2 I193 (nwayMuxOut_1n[6], inp_1d[6], nwaySelect_0n[1]);
  ND2 I194 (nwayMuxOut_1n[7], inp_1d[7], nwaySelect_0n[1]);
  ND2 I195 (nwayMuxOut_1n[8], inp_1d[8], nwaySelect_0n[1]);
  ND2 I196 (nwayMuxOut_1n[9], inp_1d[9], nwaySelect_0n[1]);
  ND2 I197 (nwayMuxOut_1n[10], inp_1d[10], nwaySelect_0n[1]);
  ND2 I198 (nwayMuxOut_1n[11], inp_1d[11], nwaySelect_0n[1]);
  ND2 I199 (nwayMuxOut_1n[12], inp_1d[12], nwaySelect_0n[1]);
  ND2 I200 (nwayMuxOut_1n[13], inp_1d[13], nwaySelect_0n[1]);
  ND2 I201 (nwayMuxOut_1n[14], inp_1d[14], nwaySelect_0n[1]);
  ND2 I202 (nwayMuxOut_1n[15], inp_1d[15], nwaySelect_0n[1]);
  ND2 I203 (nwayMuxOut_1n[16], inp_1d[16], nwaySelect_0n[1]);
  ND2 I204 (nwayMuxOut_2n[0], inp_2d[0], nwaySelect_0n[2]);
  ND2 I205 (nwayMuxOut_2n[1], inp_2d[1], nwaySelect_0n[2]);
  ND2 I206 (nwayMuxOut_2n[2], inp_2d[2], nwaySelect_0n[2]);
  ND2 I207 (nwayMuxOut_2n[3], inp_2d[3], nwaySelect_0n[2]);
  ND2 I208 (nwayMuxOut_2n[4], inp_2d[4], nwaySelect_0n[2]);
  ND2 I209 (nwayMuxOut_2n[5], inp_2d[5], nwaySelect_0n[2]);
  ND2 I210 (nwayMuxOut_2n[6], inp_2d[6], nwaySelect_0n[2]);
  ND2 I211 (nwayMuxOut_2n[7], inp_2d[7], nwaySelect_0n[2]);
  ND2 I212 (nwayMuxOut_2n[8], inp_2d[8], nwaySelect_0n[2]);
  ND2 I213 (nwayMuxOut_2n[9], inp_2d[9], nwaySelect_0n[2]);
  ND2 I214 (nwayMuxOut_2n[10], inp_2d[10], nwaySelect_0n[2]);
  ND2 I215 (nwayMuxOut_2n[11], inp_2d[11], nwaySelect_0n[2]);
  ND2 I216 (nwayMuxOut_2n[12], inp_2d[12], nwaySelect_0n[2]);
  ND2 I217 (nwayMuxOut_2n[13], inp_2d[13], nwaySelect_0n[2]);
  ND2 I218 (nwayMuxOut_2n[14], inp_2d[14], nwaySelect_0n[2]);
  ND2 I219 (nwayMuxOut_2n[15], inp_2d[15], nwaySelect_0n[2]);
  ND2 I220 (nwayMuxOut_2n[16], inp_2d[16], nwaySelect_0n[2]);
  ND2 I221 (nwayMuxOut_3n[0], inp_3d[0], nwaySelect_0n[3]);
  ND2 I222 (nwayMuxOut_3n[1], inp_3d[1], nwaySelect_0n[3]);
  ND2 I223 (nwayMuxOut_3n[2], inp_3d[2], nwaySelect_0n[3]);
  ND2 I224 (nwayMuxOut_3n[3], inp_3d[3], nwaySelect_0n[3]);
  ND2 I225 (nwayMuxOut_3n[4], inp_3d[4], nwaySelect_0n[3]);
  ND2 I226 (nwayMuxOut_3n[5], inp_3d[5], nwaySelect_0n[3]);
  ND2 I227 (nwayMuxOut_3n[6], inp_3d[6], nwaySelect_0n[3]);
  ND2 I228 (nwayMuxOut_3n[7], inp_3d[7], nwaySelect_0n[3]);
  ND2 I229 (nwayMuxOut_3n[8], inp_3d[8], nwaySelect_0n[3]);
  ND2 I230 (nwayMuxOut_3n[9], inp_3d[9], nwaySelect_0n[3]);
  ND2 I231 (nwayMuxOut_3n[10], inp_3d[10], nwaySelect_0n[3]);
  ND2 I232 (nwayMuxOut_3n[11], inp_3d[11], nwaySelect_0n[3]);
  ND2 I233 (nwayMuxOut_3n[12], inp_3d[12], nwaySelect_0n[3]);
  ND2 I234 (nwayMuxOut_3n[13], inp_3d[13], nwaySelect_0n[3]);
  ND2 I235 (nwayMuxOut_3n[14], inp_3d[14], nwaySelect_0n[3]);
  ND2 I236 (nwayMuxOut_3n[15], inp_3d[15], nwaySelect_0n[3]);
  ND2 I237 (nwayMuxOut_3n[16], inp_3d[16], nwaySelect_0n[3]);
  ND2 I238 (nwayMuxOut_4n[0], inp_4d[0], nwaySelect_0n[4]);
  ND2 I239 (nwayMuxOut_4n[1], inp_4d[1], nwaySelect_0n[4]);
  ND2 I240 (nwayMuxOut_4n[2], inp_4d[2], nwaySelect_0n[4]);
  ND2 I241 (nwayMuxOut_4n[3], inp_4d[3], nwaySelect_0n[4]);
  ND2 I242 (nwayMuxOut_4n[4], inp_4d[4], nwaySelect_0n[4]);
  ND2 I243 (nwayMuxOut_4n[5], inp_4d[5], nwaySelect_0n[4]);
  ND2 I244 (nwayMuxOut_4n[6], inp_4d[6], nwaySelect_0n[4]);
  ND2 I245 (nwayMuxOut_4n[7], inp_4d[7], nwaySelect_0n[4]);
  ND2 I246 (nwayMuxOut_4n[8], inp_4d[8], nwaySelect_0n[4]);
  ND2 I247 (nwayMuxOut_4n[9], inp_4d[9], nwaySelect_0n[4]);
  ND2 I248 (nwayMuxOut_4n[10], inp_4d[10], nwaySelect_0n[4]);
  ND2 I249 (nwayMuxOut_4n[11], inp_4d[11], nwaySelect_0n[4]);
  ND2 I250 (nwayMuxOut_4n[12], inp_4d[12], nwaySelect_0n[4]);
  ND2 I251 (nwayMuxOut_4n[13], inp_4d[13], nwaySelect_0n[4]);
  ND2 I252 (nwayMuxOut_4n[14], inp_4d[14], nwaySelect_0n[4]);
  ND2 I253 (nwayMuxOut_4n[15], inp_4d[15], nwaySelect_0n[4]);
  ND2 I254 (nwayMuxOut_4n[16], inp_4d[16], nwaySelect_0n[4]);
  ND2 I255 (nwayMuxOut_5n[0], inp_5d[0], nwaySelect_0n[5]);
  ND2 I256 (nwayMuxOut_5n[1], inp_5d[1], nwaySelect_0n[5]);
  ND2 I257 (nwayMuxOut_5n[2], inp_5d[2], nwaySelect_0n[5]);
  ND2 I258 (nwayMuxOut_5n[3], inp_5d[3], nwaySelect_0n[5]);
  ND2 I259 (nwayMuxOut_5n[4], inp_5d[4], nwaySelect_0n[5]);
  ND2 I260 (nwayMuxOut_5n[5], inp_5d[5], nwaySelect_0n[5]);
  ND2 I261 (nwayMuxOut_5n[6], inp_5d[6], nwaySelect_0n[5]);
  ND2 I262 (nwayMuxOut_5n[7], inp_5d[7], nwaySelect_0n[5]);
  ND2 I263 (nwayMuxOut_5n[8], inp_5d[8], nwaySelect_0n[5]);
  ND2 I264 (nwayMuxOut_5n[9], inp_5d[9], nwaySelect_0n[5]);
  ND2 I265 (nwayMuxOut_5n[10], inp_5d[10], nwaySelect_0n[5]);
  ND2 I266 (nwayMuxOut_5n[11], inp_5d[11], nwaySelect_0n[5]);
  ND2 I267 (nwayMuxOut_5n[12], inp_5d[12], nwaySelect_0n[5]);
  ND2 I268 (nwayMuxOut_5n[13], inp_5d[13], nwaySelect_0n[5]);
  ND2 I269 (nwayMuxOut_5n[14], inp_5d[14], nwaySelect_0n[5]);
  ND2 I270 (nwayMuxOut_5n[15], inp_5d[15], nwaySelect_0n[5]);
  ND2 I271 (nwayMuxOut_5n[16], inp_5d[16], nwaySelect_0n[5]);
  ND2 I272 (nwayMuxOut_6n[0], inp_6d[0], nwaySelect_0n[6]);
  ND2 I273 (nwayMuxOut_6n[1], inp_6d[1], nwaySelect_0n[6]);
  ND2 I274 (nwayMuxOut_6n[2], inp_6d[2], nwaySelect_0n[6]);
  ND2 I275 (nwayMuxOut_6n[3], inp_6d[3], nwaySelect_0n[6]);
  ND2 I276 (nwayMuxOut_6n[4], inp_6d[4], nwaySelect_0n[6]);
  ND2 I277 (nwayMuxOut_6n[5], inp_6d[5], nwaySelect_0n[6]);
  ND2 I278 (nwayMuxOut_6n[6], inp_6d[6], nwaySelect_0n[6]);
  ND2 I279 (nwayMuxOut_6n[7], inp_6d[7], nwaySelect_0n[6]);
  ND2 I280 (nwayMuxOut_6n[8], inp_6d[8], nwaySelect_0n[6]);
  ND2 I281 (nwayMuxOut_6n[9], inp_6d[9], nwaySelect_0n[6]);
  ND2 I282 (nwayMuxOut_6n[10], inp_6d[10], nwaySelect_0n[6]);
  ND2 I283 (nwayMuxOut_6n[11], inp_6d[11], nwaySelect_0n[6]);
  ND2 I284 (nwayMuxOut_6n[12], inp_6d[12], nwaySelect_0n[6]);
  ND2 I285 (nwayMuxOut_6n[13], inp_6d[13], nwaySelect_0n[6]);
  ND2 I286 (nwayMuxOut_6n[14], inp_6d[14], nwaySelect_0n[6]);
  ND2 I287 (nwayMuxOut_6n[15], inp_6d[15], nwaySelect_0n[6]);
  ND2 I288 (nwayMuxOut_6n[16], inp_6d[16], nwaySelect_0n[6]);
  ND2 I289 (nwayMuxOut_7n[0], inp_7d[0], nwaySelect_0n[7]);
  ND2 I290 (nwayMuxOut_7n[1], inp_7d[1], nwaySelect_0n[7]);
  ND2 I291 (nwayMuxOut_7n[2], inp_7d[2], nwaySelect_0n[7]);
  ND2 I292 (nwayMuxOut_7n[3], inp_7d[3], nwaySelect_0n[7]);
  ND2 I293 (nwayMuxOut_7n[4], inp_7d[4], nwaySelect_0n[7]);
  ND2 I294 (nwayMuxOut_7n[5], inp_7d[5], nwaySelect_0n[7]);
  ND2 I295 (nwayMuxOut_7n[6], inp_7d[6], nwaySelect_0n[7]);
  ND2 I296 (nwayMuxOut_7n[7], inp_7d[7], nwaySelect_0n[7]);
  ND2 I297 (nwayMuxOut_7n[8], inp_7d[8], nwaySelect_0n[7]);
  ND2 I298 (nwayMuxOut_7n[9], inp_7d[9], nwaySelect_0n[7]);
  ND2 I299 (nwayMuxOut_7n[10], inp_7d[10], nwaySelect_0n[7]);
  ND2 I300 (nwayMuxOut_7n[11], inp_7d[11], nwaySelect_0n[7]);
  ND2 I301 (nwayMuxOut_7n[12], inp_7d[12], nwaySelect_0n[7]);
  ND2 I302 (nwayMuxOut_7n[13], inp_7d[13], nwaySelect_0n[7]);
  ND2 I303 (nwayMuxOut_7n[14], inp_7d[14], nwaySelect_0n[7]);
  ND2 I304 (nwayMuxOut_7n[15], inp_7d[15], nwaySelect_0n[7]);
  ND2 I305 (nwayMuxOut_7n[16], inp_7d[16], nwaySelect_0n[7]);
  ND2 I306 (nwayMuxOut_8n[0], inp_8d[0], nwaySelect_0n[8]);
  ND2 I307 (nwayMuxOut_8n[1], inp_8d[1], nwaySelect_0n[8]);
  ND2 I308 (nwayMuxOut_8n[2], inp_8d[2], nwaySelect_0n[8]);
  ND2 I309 (nwayMuxOut_8n[3], inp_8d[3], nwaySelect_0n[8]);
  ND2 I310 (nwayMuxOut_8n[4], inp_8d[4], nwaySelect_0n[8]);
  ND2 I311 (nwayMuxOut_8n[5], inp_8d[5], nwaySelect_0n[8]);
  ND2 I312 (nwayMuxOut_8n[6], inp_8d[6], nwaySelect_0n[8]);
  ND2 I313 (nwayMuxOut_8n[7], inp_8d[7], nwaySelect_0n[8]);
  ND2 I314 (nwayMuxOut_8n[8], inp_8d[8], nwaySelect_0n[8]);
  ND2 I315 (nwayMuxOut_8n[9], inp_8d[9], nwaySelect_0n[8]);
  ND2 I316 (nwayMuxOut_8n[10], inp_8d[10], nwaySelect_0n[8]);
  ND2 I317 (nwayMuxOut_8n[11], inp_8d[11], nwaySelect_0n[8]);
  ND2 I318 (nwayMuxOut_8n[12], inp_8d[12], nwaySelect_0n[8]);
  ND2 I319 (nwayMuxOut_8n[13], inp_8d[13], nwaySelect_0n[8]);
  ND2 I320 (nwayMuxOut_8n[14], inp_8d[14], nwaySelect_0n[8]);
  ND2 I321 (nwayMuxOut_8n[15], inp_8d[15], nwaySelect_0n[8]);
  ND2 I322 (nwayMuxOut_8n[16], inp_8d[16], nwaySelect_0n[8]);
  ND2 I323 (nwayMuxOut_9n[0], inp_9d[0], nwaySelect_0n[9]);
  ND2 I324 (nwayMuxOut_9n[1], inp_9d[1], nwaySelect_0n[9]);
  ND2 I325 (nwayMuxOut_9n[2], inp_9d[2], nwaySelect_0n[9]);
  ND2 I326 (nwayMuxOut_9n[3], inp_9d[3], nwaySelect_0n[9]);
  ND2 I327 (nwayMuxOut_9n[4], inp_9d[4], nwaySelect_0n[9]);
  ND2 I328 (nwayMuxOut_9n[5], inp_9d[5], nwaySelect_0n[9]);
  ND2 I329 (nwayMuxOut_9n[6], inp_9d[6], nwaySelect_0n[9]);
  ND2 I330 (nwayMuxOut_9n[7], inp_9d[7], nwaySelect_0n[9]);
  ND2 I331 (nwayMuxOut_9n[8], inp_9d[8], nwaySelect_0n[9]);
  ND2 I332 (nwayMuxOut_9n[9], inp_9d[9], nwaySelect_0n[9]);
  ND2 I333 (nwayMuxOut_9n[10], inp_9d[10], nwaySelect_0n[9]);
  ND2 I334 (nwayMuxOut_9n[11], inp_9d[11], nwaySelect_0n[9]);
  ND2 I335 (nwayMuxOut_9n[12], inp_9d[12], nwaySelect_0n[9]);
  ND2 I336 (nwayMuxOut_9n[13], inp_9d[13], nwaySelect_0n[9]);
  ND2 I337 (nwayMuxOut_9n[14], inp_9d[14], nwaySelect_0n[9]);
  ND2 I338 (nwayMuxOut_9n[15], inp_9d[15], nwaySelect_0n[9]);
  ND2 I339 (nwayMuxOut_9n[16], inp_9d[16], nwaySelect_0n[9]);
  ND2 I340 (nwayMuxOut_10n[0], inp_10d[0], nwaySelect_0n[10]);
  ND2 I341 (nwayMuxOut_10n[1], inp_10d[1], nwaySelect_0n[10]);
  ND2 I342 (nwayMuxOut_10n[2], inp_10d[2], nwaySelect_0n[10]);
  ND2 I343 (nwayMuxOut_10n[3], inp_10d[3], nwaySelect_0n[10]);
  ND2 I344 (nwayMuxOut_10n[4], inp_10d[4], nwaySelect_0n[10]);
  ND2 I345 (nwayMuxOut_10n[5], inp_10d[5], nwaySelect_0n[10]);
  ND2 I346 (nwayMuxOut_10n[6], inp_10d[6], nwaySelect_0n[10]);
  ND2 I347 (nwayMuxOut_10n[7], inp_10d[7], nwaySelect_0n[10]);
  ND2 I348 (nwayMuxOut_10n[8], inp_10d[8], nwaySelect_0n[10]);
  ND2 I349 (nwayMuxOut_10n[9], inp_10d[9], nwaySelect_0n[10]);
  ND2 I350 (nwayMuxOut_10n[10], inp_10d[10], nwaySelect_0n[10]);
  ND2 I351 (nwayMuxOut_10n[11], inp_10d[11], nwaySelect_0n[10]);
  ND2 I352 (nwayMuxOut_10n[12], inp_10d[12], nwaySelect_0n[10]);
  ND2 I353 (nwayMuxOut_10n[13], inp_10d[13], nwaySelect_0n[10]);
  ND2 I354 (nwayMuxOut_10n[14], inp_10d[14], nwaySelect_0n[10]);
  ND2 I355 (nwayMuxOut_10n[15], inp_10d[15], nwaySelect_0n[10]);
  ND2 I356 (nwayMuxOut_10n[16], inp_10d[16], nwaySelect_0n[10]);
  ND2 I357 (nwayMuxOut_11n[0], inp_11d[0], nwaySelect_0n[11]);
  ND2 I358 (nwayMuxOut_11n[1], inp_11d[1], nwaySelect_0n[11]);
  ND2 I359 (nwayMuxOut_11n[2], inp_11d[2], nwaySelect_0n[11]);
  ND2 I360 (nwayMuxOut_11n[3], inp_11d[3], nwaySelect_0n[11]);
  ND2 I361 (nwayMuxOut_11n[4], inp_11d[4], nwaySelect_0n[11]);
  ND2 I362 (nwayMuxOut_11n[5], inp_11d[5], nwaySelect_0n[11]);
  ND2 I363 (nwayMuxOut_11n[6], inp_11d[6], nwaySelect_0n[11]);
  ND2 I364 (nwayMuxOut_11n[7], inp_11d[7], nwaySelect_0n[11]);
  ND2 I365 (nwayMuxOut_11n[8], inp_11d[8], nwaySelect_0n[11]);
  ND2 I366 (nwayMuxOut_11n[9], inp_11d[9], nwaySelect_0n[11]);
  ND2 I367 (nwayMuxOut_11n[10], inp_11d[10], nwaySelect_0n[11]);
  ND2 I368 (nwayMuxOut_11n[11], inp_11d[11], nwaySelect_0n[11]);
  ND2 I369 (nwayMuxOut_11n[12], inp_11d[12], nwaySelect_0n[11]);
  ND2 I370 (nwayMuxOut_11n[13], inp_11d[13], nwaySelect_0n[11]);
  ND2 I371 (nwayMuxOut_11n[14], inp_11d[14], nwaySelect_0n[11]);
  ND2 I372 (nwayMuxOut_11n[15], inp_11d[15], nwaySelect_0n[11]);
  ND2 I373 (nwayMuxOut_11n[16], inp_11d[16], nwaySelect_0n[11]);
  ND2 I374 (nwayMuxOut_12n[0], inp_12d[0], nwaySelect_0n[12]);
  ND2 I375 (nwayMuxOut_12n[1], inp_12d[1], nwaySelect_0n[12]);
  ND2 I376 (nwayMuxOut_12n[2], inp_12d[2], nwaySelect_0n[12]);
  ND2 I377 (nwayMuxOut_12n[3], inp_12d[3], nwaySelect_0n[12]);
  ND2 I378 (nwayMuxOut_12n[4], inp_12d[4], nwaySelect_0n[12]);
  ND2 I379 (nwayMuxOut_12n[5], inp_12d[5], nwaySelect_0n[12]);
  ND2 I380 (nwayMuxOut_12n[6], inp_12d[6], nwaySelect_0n[12]);
  ND2 I381 (nwayMuxOut_12n[7], inp_12d[7], nwaySelect_0n[12]);
  ND2 I382 (nwayMuxOut_12n[8], inp_12d[8], nwaySelect_0n[12]);
  ND2 I383 (nwayMuxOut_12n[9], inp_12d[9], nwaySelect_0n[12]);
  ND2 I384 (nwayMuxOut_12n[10], inp_12d[10], nwaySelect_0n[12]);
  ND2 I385 (nwayMuxOut_12n[11], inp_12d[11], nwaySelect_0n[12]);
  ND2 I386 (nwayMuxOut_12n[12], inp_12d[12], nwaySelect_0n[12]);
  ND2 I387 (nwayMuxOut_12n[13], inp_12d[13], nwaySelect_0n[12]);
  ND2 I388 (nwayMuxOut_12n[14], inp_12d[14], nwaySelect_0n[12]);
  ND2 I389 (nwayMuxOut_12n[15], inp_12d[15], nwaySelect_0n[12]);
  ND2 I390 (nwayMuxOut_12n[16], inp_12d[16], nwaySelect_0n[12]);
  ND2 I391 (nwayMuxOut_13n[0], inp_13d[0], nwaySelect_0n[13]);
  ND2 I392 (nwayMuxOut_13n[1], inp_13d[1], nwaySelect_0n[13]);
  ND2 I393 (nwayMuxOut_13n[2], inp_13d[2], nwaySelect_0n[13]);
  ND2 I394 (nwayMuxOut_13n[3], inp_13d[3], nwaySelect_0n[13]);
  ND2 I395 (nwayMuxOut_13n[4], inp_13d[4], nwaySelect_0n[13]);
  ND2 I396 (nwayMuxOut_13n[5], inp_13d[5], nwaySelect_0n[13]);
  ND2 I397 (nwayMuxOut_13n[6], inp_13d[6], nwaySelect_0n[13]);
  ND2 I398 (nwayMuxOut_13n[7], inp_13d[7], nwaySelect_0n[13]);
  ND2 I399 (nwayMuxOut_13n[8], inp_13d[8], nwaySelect_0n[13]);
  ND2 I400 (nwayMuxOut_13n[9], inp_13d[9], nwaySelect_0n[13]);
  ND2 I401 (nwayMuxOut_13n[10], inp_13d[10], nwaySelect_0n[13]);
  ND2 I402 (nwayMuxOut_13n[11], inp_13d[11], nwaySelect_0n[13]);
  ND2 I403 (nwayMuxOut_13n[12], inp_13d[12], nwaySelect_0n[13]);
  ND2 I404 (nwayMuxOut_13n[13], inp_13d[13], nwaySelect_0n[13]);
  ND2 I405 (nwayMuxOut_13n[14], inp_13d[14], nwaySelect_0n[13]);
  ND2 I406 (nwayMuxOut_13n[15], inp_13d[15], nwaySelect_0n[13]);
  ND2 I407 (nwayMuxOut_13n[16], inp_13d[16], nwaySelect_0n[13]);
  ND2 I408 (nwayMuxOut_14n[0], inp_14d[0], nwaySelect_0n[14]);
  ND2 I409 (nwayMuxOut_14n[1], inp_14d[1], nwaySelect_0n[14]);
  ND2 I410 (nwayMuxOut_14n[2], inp_14d[2], nwaySelect_0n[14]);
  ND2 I411 (nwayMuxOut_14n[3], inp_14d[3], nwaySelect_0n[14]);
  ND2 I412 (nwayMuxOut_14n[4], inp_14d[4], nwaySelect_0n[14]);
  ND2 I413 (nwayMuxOut_14n[5], inp_14d[5], nwaySelect_0n[14]);
  ND2 I414 (nwayMuxOut_14n[6], inp_14d[6], nwaySelect_0n[14]);
  ND2 I415 (nwayMuxOut_14n[7], inp_14d[7], nwaySelect_0n[14]);
  ND2 I416 (nwayMuxOut_14n[8], inp_14d[8], nwaySelect_0n[14]);
  ND2 I417 (nwayMuxOut_14n[9], inp_14d[9], nwaySelect_0n[14]);
  ND2 I418 (nwayMuxOut_14n[10], inp_14d[10], nwaySelect_0n[14]);
  ND2 I419 (nwayMuxOut_14n[11], inp_14d[11], nwaySelect_0n[14]);
  ND2 I420 (nwayMuxOut_14n[12], inp_14d[12], nwaySelect_0n[14]);
  ND2 I421 (nwayMuxOut_14n[13], inp_14d[13], nwaySelect_0n[14]);
  ND2 I422 (nwayMuxOut_14n[14], inp_14d[14], nwaySelect_0n[14]);
  ND2 I423 (nwayMuxOut_14n[15], inp_14d[15], nwaySelect_0n[14]);
  ND2 I424 (nwayMuxOut_14n[16], inp_14d[16], nwaySelect_0n[14]);
  ND2 I425 (nwayMuxOut_15n[0], inp_15d[0], nwaySelect_0n[15]);
  ND2 I426 (nwayMuxOut_15n[1], inp_15d[1], nwaySelect_0n[15]);
  ND2 I427 (nwayMuxOut_15n[2], inp_15d[2], nwaySelect_0n[15]);
  ND2 I428 (nwayMuxOut_15n[3], inp_15d[3], nwaySelect_0n[15]);
  ND2 I429 (nwayMuxOut_15n[4], inp_15d[4], nwaySelect_0n[15]);
  ND2 I430 (nwayMuxOut_15n[5], inp_15d[5], nwaySelect_0n[15]);
  ND2 I431 (nwayMuxOut_15n[6], inp_15d[6], nwaySelect_0n[15]);
  ND2 I432 (nwayMuxOut_15n[7], inp_15d[7], nwaySelect_0n[15]);
  ND2 I433 (nwayMuxOut_15n[8], inp_15d[8], nwaySelect_0n[15]);
  ND2 I434 (nwayMuxOut_15n[9], inp_15d[9], nwaySelect_0n[15]);
  ND2 I435 (nwayMuxOut_15n[10], inp_15d[10], nwaySelect_0n[15]);
  ND2 I436 (nwayMuxOut_15n[11], inp_15d[11], nwaySelect_0n[15]);
  ND2 I437 (nwayMuxOut_15n[12], inp_15d[12], nwaySelect_0n[15]);
  ND2 I438 (nwayMuxOut_15n[13], inp_15d[13], nwaySelect_0n[15]);
  ND2 I439 (nwayMuxOut_15n[14], inp_15d[14], nwaySelect_0n[15]);
  ND2 I440 (nwayMuxOut_15n[15], inp_15d[15], nwaySelect_0n[15]);
  ND2 I441 (nwayMuxOut_15n[16], inp_15d[16], nwaySelect_0n[15]);
  ND2 I442 (nwayMuxOut_16n[0], inp_16d[0], nwaySelect_0n[16]);
  ND2 I443 (nwayMuxOut_16n[1], inp_16d[1], nwaySelect_0n[16]);
  ND2 I444 (nwayMuxOut_16n[2], inp_16d[2], nwaySelect_0n[16]);
  ND2 I445 (nwayMuxOut_16n[3], inp_16d[3], nwaySelect_0n[16]);
  ND2 I446 (nwayMuxOut_16n[4], inp_16d[4], nwaySelect_0n[16]);
  ND2 I447 (nwayMuxOut_16n[5], inp_16d[5], nwaySelect_0n[16]);
  ND2 I448 (nwayMuxOut_16n[6], inp_16d[6], nwaySelect_0n[16]);
  ND2 I449 (nwayMuxOut_16n[7], inp_16d[7], nwaySelect_0n[16]);
  ND2 I450 (nwayMuxOut_16n[8], inp_16d[8], nwaySelect_0n[16]);
  ND2 I451 (nwayMuxOut_16n[9], inp_16d[9], nwaySelect_0n[16]);
  ND2 I452 (nwayMuxOut_16n[10], inp_16d[10], nwaySelect_0n[16]);
  ND2 I453 (nwayMuxOut_16n[11], inp_16d[11], nwaySelect_0n[16]);
  ND2 I454 (nwayMuxOut_16n[12], inp_16d[12], nwaySelect_0n[16]);
  ND2 I455 (nwayMuxOut_16n[13], inp_16d[13], nwaySelect_0n[16]);
  ND2 I456 (nwayMuxOut_16n[14], inp_16d[14], nwaySelect_0n[16]);
  ND2 I457 (nwayMuxOut_16n[15], inp_16d[15], nwaySelect_0n[16]);
  ND2 I458 (nwayMuxOut_16n[16], inp_16d[16], nwaySelect_0n[16]);
  ND2 I459 (nwayMuxOut_17n[0], inp_17d[0], nwaySelect_0n[17]);
  ND2 I460 (nwayMuxOut_17n[1], inp_17d[1], nwaySelect_0n[17]);
  ND2 I461 (nwayMuxOut_17n[2], inp_17d[2], nwaySelect_0n[17]);
  ND2 I462 (nwayMuxOut_17n[3], inp_17d[3], nwaySelect_0n[17]);
  ND2 I463 (nwayMuxOut_17n[4], inp_17d[4], nwaySelect_0n[17]);
  ND2 I464 (nwayMuxOut_17n[5], inp_17d[5], nwaySelect_0n[17]);
  ND2 I465 (nwayMuxOut_17n[6], inp_17d[6], nwaySelect_0n[17]);
  ND2 I466 (nwayMuxOut_17n[7], inp_17d[7], nwaySelect_0n[17]);
  ND2 I467 (nwayMuxOut_17n[8], inp_17d[8], nwaySelect_0n[17]);
  ND2 I468 (nwayMuxOut_17n[9], inp_17d[9], nwaySelect_0n[17]);
  ND2 I469 (nwayMuxOut_17n[10], inp_17d[10], nwaySelect_0n[17]);
  ND2 I470 (nwayMuxOut_17n[11], inp_17d[11], nwaySelect_0n[17]);
  ND2 I471 (nwayMuxOut_17n[12], inp_17d[12], nwaySelect_0n[17]);
  ND2 I472 (nwayMuxOut_17n[13], inp_17d[13], nwaySelect_0n[17]);
  ND2 I473 (nwayMuxOut_17n[14], inp_17d[14], nwaySelect_0n[17]);
  ND2 I474 (nwayMuxOut_17n[15], inp_17d[15], nwaySelect_0n[17]);
  ND2 I475 (nwayMuxOut_17n[16], inp_17d[16], nwaySelect_0n[17]);
  ND2 I476 (nwayMuxOut_18n[0], inp_18d[0], nwaySelect_0n[18]);
  ND2 I477 (nwayMuxOut_18n[1], inp_18d[1], nwaySelect_0n[18]);
  ND2 I478 (nwayMuxOut_18n[2], inp_18d[2], nwaySelect_0n[18]);
  ND2 I479 (nwayMuxOut_18n[3], inp_18d[3], nwaySelect_0n[18]);
  ND2 I480 (nwayMuxOut_18n[4], inp_18d[4], nwaySelect_0n[18]);
  ND2 I481 (nwayMuxOut_18n[5], inp_18d[5], nwaySelect_0n[18]);
  ND2 I482 (nwayMuxOut_18n[6], inp_18d[6], nwaySelect_0n[18]);
  ND2 I483 (nwayMuxOut_18n[7], inp_18d[7], nwaySelect_0n[18]);
  ND2 I484 (nwayMuxOut_18n[8], inp_18d[8], nwaySelect_0n[18]);
  ND2 I485 (nwayMuxOut_18n[9], inp_18d[9], nwaySelect_0n[18]);
  ND2 I486 (nwayMuxOut_18n[10], inp_18d[10], nwaySelect_0n[18]);
  ND2 I487 (nwayMuxOut_18n[11], inp_18d[11], nwaySelect_0n[18]);
  ND2 I488 (nwayMuxOut_18n[12], inp_18d[12], nwaySelect_0n[18]);
  ND2 I489 (nwayMuxOut_18n[13], inp_18d[13], nwaySelect_0n[18]);
  ND2 I490 (nwayMuxOut_18n[14], inp_18d[14], nwaySelect_0n[18]);
  ND2 I491 (nwayMuxOut_18n[15], inp_18d[15], nwaySelect_0n[18]);
  ND2 I492 (nwayMuxOut_18n[16], inp_18d[16], nwaySelect_0n[18]);
  ND2 I493 (nwayMuxOut_19n[0], inp_19d[0], nwaySelect_0n[19]);
  ND2 I494 (nwayMuxOut_19n[1], inp_19d[1], nwaySelect_0n[19]);
  ND2 I495 (nwayMuxOut_19n[2], inp_19d[2], nwaySelect_0n[19]);
  ND2 I496 (nwayMuxOut_19n[3], inp_19d[3], nwaySelect_0n[19]);
  ND2 I497 (nwayMuxOut_19n[4], inp_19d[4], nwaySelect_0n[19]);
  ND2 I498 (nwayMuxOut_19n[5], inp_19d[5], nwaySelect_0n[19]);
  ND2 I499 (nwayMuxOut_19n[6], inp_19d[6], nwaySelect_0n[19]);
  ND2 I500 (nwayMuxOut_19n[7], inp_19d[7], nwaySelect_0n[19]);
  ND2 I501 (nwayMuxOut_19n[8], inp_19d[8], nwaySelect_0n[19]);
  ND2 I502 (nwayMuxOut_19n[9], inp_19d[9], nwaySelect_0n[19]);
  ND2 I503 (nwayMuxOut_19n[10], inp_19d[10], nwaySelect_0n[19]);
  ND2 I504 (nwayMuxOut_19n[11], inp_19d[11], nwaySelect_0n[19]);
  ND2 I505 (nwayMuxOut_19n[12], inp_19d[12], nwaySelect_0n[19]);
  ND2 I506 (nwayMuxOut_19n[13], inp_19d[13], nwaySelect_0n[19]);
  ND2 I507 (nwayMuxOut_19n[14], inp_19d[14], nwaySelect_0n[19]);
  ND2 I508 (nwayMuxOut_19n[15], inp_19d[15], nwaySelect_0n[19]);
  ND2 I509 (nwayMuxOut_19n[16], inp_19d[16], nwaySelect_0n[19]);
  ND2 I510 (nwayMuxOut_20n[0], inp_20d[0], nwaySelect_0n[20]);
  ND2 I511 (nwayMuxOut_20n[1], inp_20d[1], nwaySelect_0n[20]);
  ND2 I512 (nwayMuxOut_20n[2], inp_20d[2], nwaySelect_0n[20]);
  ND2 I513 (nwayMuxOut_20n[3], inp_20d[3], nwaySelect_0n[20]);
  ND2 I514 (nwayMuxOut_20n[4], inp_20d[4], nwaySelect_0n[20]);
  ND2 I515 (nwayMuxOut_20n[5], inp_20d[5], nwaySelect_0n[20]);
  ND2 I516 (nwayMuxOut_20n[6], inp_20d[6], nwaySelect_0n[20]);
  ND2 I517 (nwayMuxOut_20n[7], inp_20d[7], nwaySelect_0n[20]);
  ND2 I518 (nwayMuxOut_20n[8], inp_20d[8], nwaySelect_0n[20]);
  ND2 I519 (nwayMuxOut_20n[9], inp_20d[9], nwaySelect_0n[20]);
  ND2 I520 (nwayMuxOut_20n[10], inp_20d[10], nwaySelect_0n[20]);
  ND2 I521 (nwayMuxOut_20n[11], inp_20d[11], nwaySelect_0n[20]);
  ND2 I522 (nwayMuxOut_20n[12], inp_20d[12], nwaySelect_0n[20]);
  ND2 I523 (nwayMuxOut_20n[13], inp_20d[13], nwaySelect_0n[20]);
  ND2 I524 (nwayMuxOut_20n[14], inp_20d[14], nwaySelect_0n[20]);
  ND2 I525 (nwayMuxOut_20n[15], inp_20d[15], nwaySelect_0n[20]);
  ND2 I526 (nwayMuxOut_20n[16], inp_20d[16], nwaySelect_0n[20]);
  ND2 I527 (nwayMuxOut_21n[0], inp_21d[0], nwaySelect_0n[21]);
  ND2 I528 (nwayMuxOut_21n[1], inp_21d[1], nwaySelect_0n[21]);
  ND2 I529 (nwayMuxOut_21n[2], inp_21d[2], nwaySelect_0n[21]);
  ND2 I530 (nwayMuxOut_21n[3], inp_21d[3], nwaySelect_0n[21]);
  ND2 I531 (nwayMuxOut_21n[4], inp_21d[4], nwaySelect_0n[21]);
  ND2 I532 (nwayMuxOut_21n[5], inp_21d[5], nwaySelect_0n[21]);
  ND2 I533 (nwayMuxOut_21n[6], inp_21d[6], nwaySelect_0n[21]);
  ND2 I534 (nwayMuxOut_21n[7], inp_21d[7], nwaySelect_0n[21]);
  ND2 I535 (nwayMuxOut_21n[8], inp_21d[8], nwaySelect_0n[21]);
  ND2 I536 (nwayMuxOut_21n[9], inp_21d[9], nwaySelect_0n[21]);
  ND2 I537 (nwayMuxOut_21n[10], inp_21d[10], nwaySelect_0n[21]);
  ND2 I538 (nwayMuxOut_21n[11], inp_21d[11], nwaySelect_0n[21]);
  ND2 I539 (nwayMuxOut_21n[12], inp_21d[12], nwaySelect_0n[21]);
  ND2 I540 (nwayMuxOut_21n[13], inp_21d[13], nwaySelect_0n[21]);
  ND2 I541 (nwayMuxOut_21n[14], inp_21d[14], nwaySelect_0n[21]);
  ND2 I542 (nwayMuxOut_21n[15], inp_21d[15], nwaySelect_0n[21]);
  ND2 I543 (nwayMuxOut_21n[16], inp_21d[16], nwaySelect_0n[21]);
  ND2 I544 (nwayMuxOut_22n[0], inp_22d[0], nwaySelect_0n[22]);
  ND2 I545 (nwayMuxOut_22n[1], inp_22d[1], nwaySelect_0n[22]);
  ND2 I546 (nwayMuxOut_22n[2], inp_22d[2], nwaySelect_0n[22]);
  ND2 I547 (nwayMuxOut_22n[3], inp_22d[3], nwaySelect_0n[22]);
  ND2 I548 (nwayMuxOut_22n[4], inp_22d[4], nwaySelect_0n[22]);
  ND2 I549 (nwayMuxOut_22n[5], inp_22d[5], nwaySelect_0n[22]);
  ND2 I550 (nwayMuxOut_22n[6], inp_22d[6], nwaySelect_0n[22]);
  ND2 I551 (nwayMuxOut_22n[7], inp_22d[7], nwaySelect_0n[22]);
  ND2 I552 (nwayMuxOut_22n[8], inp_22d[8], nwaySelect_0n[22]);
  ND2 I553 (nwayMuxOut_22n[9], inp_22d[9], nwaySelect_0n[22]);
  ND2 I554 (nwayMuxOut_22n[10], inp_22d[10], nwaySelect_0n[22]);
  ND2 I555 (nwayMuxOut_22n[11], inp_22d[11], nwaySelect_0n[22]);
  ND2 I556 (nwayMuxOut_22n[12], inp_22d[12], nwaySelect_0n[22]);
  ND2 I557 (nwayMuxOut_22n[13], inp_22d[13], nwaySelect_0n[22]);
  ND2 I558 (nwayMuxOut_22n[14], inp_22d[14], nwaySelect_0n[22]);
  ND2 I559 (nwayMuxOut_22n[15], inp_22d[15], nwaySelect_0n[22]);
  ND2 I560 (nwayMuxOut_22n[16], inp_22d[16], nwaySelect_0n[22]);
  ND2 I561 (nwayMuxOut_23n[0], inp_23d[0], nwaySelect_0n[23]);
  ND2 I562 (nwayMuxOut_23n[1], inp_23d[1], nwaySelect_0n[23]);
  ND2 I563 (nwayMuxOut_23n[2], inp_23d[2], nwaySelect_0n[23]);
  ND2 I564 (nwayMuxOut_23n[3], inp_23d[3], nwaySelect_0n[23]);
  ND2 I565 (nwayMuxOut_23n[4], inp_23d[4], nwaySelect_0n[23]);
  ND2 I566 (nwayMuxOut_23n[5], inp_23d[5], nwaySelect_0n[23]);
  ND2 I567 (nwayMuxOut_23n[6], inp_23d[6], nwaySelect_0n[23]);
  ND2 I568 (nwayMuxOut_23n[7], inp_23d[7], nwaySelect_0n[23]);
  ND2 I569 (nwayMuxOut_23n[8], inp_23d[8], nwaySelect_0n[23]);
  ND2 I570 (nwayMuxOut_23n[9], inp_23d[9], nwaySelect_0n[23]);
  ND2 I571 (nwayMuxOut_23n[10], inp_23d[10], nwaySelect_0n[23]);
  ND2 I572 (nwayMuxOut_23n[11], inp_23d[11], nwaySelect_0n[23]);
  ND2 I573 (nwayMuxOut_23n[12], inp_23d[12], nwaySelect_0n[23]);
  ND2 I574 (nwayMuxOut_23n[13], inp_23d[13], nwaySelect_0n[23]);
  ND2 I575 (nwayMuxOut_23n[14], inp_23d[14], nwaySelect_0n[23]);
  ND2 I576 (nwayMuxOut_23n[15], inp_23d[15], nwaySelect_0n[23]);
  ND2 I577 (nwayMuxOut_23n[16], inp_23d[16], nwaySelect_0n[23]);
  ND2 I578 (nwayMuxOut_24n[0], inp_24d[0], nwaySelect_0n[24]);
  ND2 I579 (nwayMuxOut_24n[1], inp_24d[1], nwaySelect_0n[24]);
  ND2 I580 (nwayMuxOut_24n[2], inp_24d[2], nwaySelect_0n[24]);
  ND2 I581 (nwayMuxOut_24n[3], inp_24d[3], nwaySelect_0n[24]);
  ND2 I582 (nwayMuxOut_24n[4], inp_24d[4], nwaySelect_0n[24]);
  ND2 I583 (nwayMuxOut_24n[5], inp_24d[5], nwaySelect_0n[24]);
  ND2 I584 (nwayMuxOut_24n[6], inp_24d[6], nwaySelect_0n[24]);
  ND2 I585 (nwayMuxOut_24n[7], inp_24d[7], nwaySelect_0n[24]);
  ND2 I586 (nwayMuxOut_24n[8], inp_24d[8], nwaySelect_0n[24]);
  ND2 I587 (nwayMuxOut_24n[9], inp_24d[9], nwaySelect_0n[24]);
  ND2 I588 (nwayMuxOut_24n[10], inp_24d[10], nwaySelect_0n[24]);
  ND2 I589 (nwayMuxOut_24n[11], inp_24d[11], nwaySelect_0n[24]);
  ND2 I590 (nwayMuxOut_24n[12], inp_24d[12], nwaySelect_0n[24]);
  ND2 I591 (nwayMuxOut_24n[13], inp_24d[13], nwaySelect_0n[24]);
  ND2 I592 (nwayMuxOut_24n[14], inp_24d[14], nwaySelect_0n[24]);
  ND2 I593 (nwayMuxOut_24n[15], inp_24d[15], nwaySelect_0n[24]);
  ND2 I594 (nwayMuxOut_24n[16], inp_24d[16], nwaySelect_0n[24]);
  OR2 I595 (nwaySelect_0n[0], inp_0a, inp_0r);
  OR2 I596 (nwaySelect_0n[1], inp_1a, inp_1r);
  OR2 I597 (nwaySelect_0n[2], inp_2a, inp_2r);
  OR2 I598 (nwaySelect_0n[3], inp_3a, inp_3r);
  OR2 I599 (nwaySelect_0n[4], inp_4a, inp_4r);
  OR2 I600 (nwaySelect_0n[5], inp_5a, inp_5r);
  OR2 I601 (nwaySelect_0n[6], inp_6a, inp_6r);
  OR2 I602 (nwaySelect_0n[7], inp_7a, inp_7r);
  OR2 I603 (nwaySelect_0n[8], inp_8a, inp_8r);
  OR2 I604 (nwaySelect_0n[9], inp_9a, inp_9r);
  OR2 I605 (nwaySelect_0n[10], inp_10a, inp_10r);
  OR2 I606 (nwaySelect_0n[11], inp_11a, inp_11r);
  OR2 I607 (nwaySelect_0n[12], inp_12a, inp_12r);
  OR2 I608 (nwaySelect_0n[13], inp_13a, inp_13r);
  OR2 I609 (nwaySelect_0n[14], inp_14a, inp_14r);
  OR2 I610 (nwaySelect_0n[15], inp_15a, inp_15r);
  OR2 I611 (nwaySelect_0n[16], inp_16a, inp_16r);
  OR2 I612 (nwaySelect_0n[17], inp_17a, inp_17r);
  OR2 I613 (nwaySelect_0n[18], inp_18a, inp_18r);
  OR2 I614 (nwaySelect_0n[19], inp_19a, inp_19r);
  OR2 I615 (nwaySelect_0n[20], inp_20a, inp_20r);
  OR2 I616 (nwaySelect_0n[21], inp_21a, inp_21r);
  OR2 I617 (nwaySelect_0n[22], inp_22a, inp_22r);
  OR2 I618 (nwaySelect_0n[23], inp_23a, inp_23r);
  OR2 I619 (nwaySelect_0n[24], inp_24a, inp_24r);
  C2 I620 (inp_0a, inp_0r, out_0a);
  C2 I621 (inp_1a, inp_1r, out_0a);
  C2 I622 (inp_2a, inp_2r, out_0a);
  C2 I623 (inp_3a, inp_3r, out_0a);
  C2 I624 (inp_4a, inp_4r, out_0a);
  C2 I625 (inp_5a, inp_5r, out_0a);
  C2 I626 (inp_6a, inp_6r, out_0a);
  C2 I627 (inp_7a, inp_7r, out_0a);
  C2 I628 (inp_8a, inp_8r, out_0a);
  C2 I629 (inp_9a, inp_9r, out_0a);
  C2 I630 (inp_10a, inp_10r, out_0a);
  C2 I631 (inp_11a, inp_11r, out_0a);
  C2 I632 (inp_12a, inp_12r, out_0a);
  C2 I633 (inp_13a, inp_13r, out_0a);
  C2 I634 (inp_14a, inp_14r, out_0a);
  C2 I635 (inp_15a, inp_15r, out_0a);
  C2 I636 (inp_16a, inp_16r, out_0a);
  C2 I637 (inp_17a, inp_17r, out_0a);
  C2 I638 (inp_18a, inp_18r, out_0a);
  C2 I639 (inp_19a, inp_19r, out_0a);
  C2 I640 (inp_20a, inp_20r, out_0a);
  C2 I641 (inp_21a, inp_21r, out_0a);
  C2 I642 (inp_22a, inp_22r, out_0a);
  C2 I643 (inp_23a, inp_23r, out_0a);
  C2 I644 (inp_24a, inp_24r, out_0a);
  NR4 I645 (internal_0n[153], inp_0r, inp_1r, inp_2r, inp_3r);
  NR4 I646 (internal_0n[154], inp_4r, inp_5r, inp_6r, inp_7r);
  NR4 I647 (internal_0n[155], inp_8r, inp_9r, inp_10r, inp_11r);
  NR4 I648 (internal_0n[156], inp_12r, inp_13r, inp_14r, inp_15r);
  NR4 I649 (internal_0n[157], inp_16r, inp_17r, inp_18r, inp_19r);
  NR2 I650 (internal_0n[158], inp_20r, inp_21r);
  NR3 I651 (internal_0n[159], inp_22r, inp_23r, inp_24r);
  ND4 I652 (internal_0n[160], internal_0n[153], internal_0n[154], internal_0n[155], internal_0n[156]);
  ND3 I653 (internal_0n[161], internal_0n[157], internal_0n[158], internal_0n[159]);
  OR2 I654 (out_0r, internal_0n[160], internal_0n[161]);
endmodule

module BrzCase_1_2_s5_0_3b1 (
  inp_0r, inp_0a, inp_0d,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a
);
  input inp_0r;
  output inp_0a;
  input inp_0d;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  wire t_0n;
  wire c_0n;
  wire elseAck_0n;
  wire [1:0] int0_0n;
  OR2 I0 (inp_0a, activateOut_0a, activateOut_1a);
  assign int0_0n[0] = c_0n;
  assign int0_0n[1] = t_0n;
  assign activateOut_1r = int0_0n[1];
  assign activateOut_0r = int0_0n[0];
  demux2 I5 (inp_0r, c_0n, t_0n, inp_0d);
endmodule

module BrzCombine_9_1_8 (
  out_0r, out_0a, out_0d,
  LSInp_0r, LSInp_0a, LSInp_0d,
  MSInp_0r, MSInp_0a, MSInp_0d
);
  input out_0r;
  output out_0a;
  output [8:0] out_0d;
  output LSInp_0r;
  input LSInp_0a;
  input LSInp_0d;
  output MSInp_0r;
  input MSInp_0a;
  input [7:0] MSInp_0d;
  C2 I0 (out_0a, LSInp_0a, MSInp_0a);
  assign LSInp_0r = out_0r;
  assign MSInp_0r = out_0r;
  assign out_0d[0] = LSInp_0d;
  assign out_0d[1] = MSInp_0d[0];
  assign out_0d[2] = MSInp_0d[1];
  assign out_0d[3] = MSInp_0d[2];
  assign out_0d[4] = MSInp_0d[3];
  assign out_0d[5] = MSInp_0d[4];
  assign out_0d[6] = MSInp_0d[5];
  assign out_0d[7] = MSInp_0d[6];
  assign out_0d[8] = MSInp_0d[7];
endmodule

module BrzCombine_17_9_8 (
  out_0r, out_0a, out_0d,
  LSInp_0r, LSInp_0a, LSInp_0d,
  MSInp_0r, MSInp_0a, MSInp_0d
);
  input out_0r;
  output out_0a;
  output [16:0] out_0d;
  output LSInp_0r;
  input LSInp_0a;
  input [8:0] LSInp_0d;
  output MSInp_0r;
  input MSInp_0a;
  input [7:0] MSInp_0d;
  C2 I0 (out_0a, LSInp_0a, MSInp_0a);
  assign LSInp_0r = out_0r;
  assign MSInp_0r = out_0r;
  assign out_0d[0] = LSInp_0d[0];
  assign out_0d[1] = LSInp_0d[1];
  assign out_0d[2] = LSInp_0d[2];
  assign out_0d[3] = LSInp_0d[3];
  assign out_0d[4] = LSInp_0d[4];
  assign out_0d[5] = LSInp_0d[5];
  assign out_0d[6] = LSInp_0d[6];
  assign out_0d[7] = LSInp_0d[7];
  assign out_0d[8] = LSInp_0d[8];
  assign out_0d[9] = MSInp_0d[0];
  assign out_0d[10] = MSInp_0d[1];
  assign out_0d[11] = MSInp_0d[2];
  assign out_0d[12] = MSInp_0d[3];
  assign out_0d[13] = MSInp_0d[4];
  assign out_0d[14] = MSInp_0d[5];
  assign out_0d[15] = MSInp_0d[6];
  assign out_0d[16] = MSInp_0d[7];
endmodule

module BrzCombine_17_16_1 (
  out_0r, out_0a, out_0d,
  LSInp_0r, LSInp_0a, LSInp_0d,
  MSInp_0r, MSInp_0a, MSInp_0d
);
  input out_0r;
  output out_0a;
  output [16:0] out_0d;
  output LSInp_0r;
  input LSInp_0a;
  input [15:0] LSInp_0d;
  output MSInp_0r;
  input MSInp_0a;
  input MSInp_0d;
  C2 I0 (out_0a, LSInp_0a, MSInp_0a);
  assign LSInp_0r = out_0r;
  assign MSInp_0r = out_0r;
  assign out_0d[0] = LSInp_0d[0];
  assign out_0d[1] = LSInp_0d[1];
  assign out_0d[2] = LSInp_0d[2];
  assign out_0d[3] = LSInp_0d[3];
  assign out_0d[4] = LSInp_0d[4];
  assign out_0d[5] = LSInp_0d[5];
  assign out_0d[6] = LSInp_0d[6];
  assign out_0d[7] = LSInp_0d[7];
  assign out_0d[8] = LSInp_0d[8];
  assign out_0d[9] = LSInp_0d[9];
  assign out_0d[10] = LSInp_0d[10];
  assign out_0d[11] = LSInp_0d[11];
  assign out_0d[12] = LSInp_0d[12];
  assign out_0d[13] = LSInp_0d[13];
  assign out_0d[14] = LSInp_0d[14];
  assign out_0d[15] = LSInp_0d[15];
  assign out_0d[16] = MSInp_0d;
endmodule

module telem (
  Ar,
  Aa,
  Br,
  Ba
);
  input Ar;
  output Aa;
  output Br;
  input Ba;
  wire s_0n;
  ACU0D1 I0 (Aa, Ba, Ar);
  IV I1 (s_0n, Aa);
  AN2 I2 (Br, Ar, s_0n);
endmodule

module BrzConcur_2 (
  activate_0r, activate_0a,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a
);
  input activate_0r;
  output activate_0a;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  wire [1:0] acks_0n;
  C2 I0 (activate_0a, acks_0n[0], acks_0n[1]);
  telem I1 (activate_0r, acks_0n[0], activateOut_0r, activateOut_0a);
  telem I2 (activate_0r, acks_0n[1], activateOut_1r, activateOut_1a);
endmodule

module BrzConcur_3 (
  activate_0r, activate_0a,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a,
  activateOut_2r, activateOut_2a
);
  input activate_0r;
  output activate_0a;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  output activateOut_2r;
  input activateOut_2a;
  wire [2:0] acks_0n;
  C3 I0 (activate_0a, acks_0n[0], acks_0n[1], acks_0n[2]);
  telem I1 (activate_0r, acks_0n[0], activateOut_0r, activateOut_0a);
  telem I2 (activate_0r, acks_0n[1], activateOut_1r, activateOut_1a);
  telem I3 (activate_0r, acks_0n[2], activateOut_2r, activateOut_2a);
endmodule

module BrzConstant_1_0 (
  out_0r, out_0a, out_0d
);
  input out_0r;
  output out_0a;
  output out_0d;
  wire gnd;
  GND gnd_cell_instance (gnd);
  assign out_0a = out_0r;
  assign out_0d = gnd;
endmodule

module BrzConstant_9_0 (
  out_0r, out_0a, out_0d
);
  input out_0r;
  output out_0a;
  output [8:0] out_0d;
  wire gnd;
  GND gnd_cell_instance (gnd);
  assign out_0a = out_0r;
  assign out_0d[0] = gnd;
  assign out_0d[1] = gnd;
  assign out_0d[2] = gnd;
  assign out_0d[3] = gnd;
  assign out_0d[4] = gnd;
  assign out_0d[5] = gnd;
  assign out_0d[6] = gnd;
  assign out_0d[7] = gnd;
  assign out_0d[8] = gnd;
endmodule

module BrzFetch_1_s5_false (
  activate_0r, activate_0a,
  inp_0r, inp_0a, inp_0d,
  out_0r, out_0a, out_0d
);
  input activate_0r;
  output activate_0a;
  output inp_0r;
  input inp_0a;
  input inp_0d;
  output out_0r;
  input out_0a;
  output out_0d;
  assign activate_0a = out_0a;
  assign out_0r = inp_0a;
  assign inp_0r = activate_0r;
  assign out_0d = inp_0d;
endmodule

module BrzFetch_8_s5_false (
  activate_0r, activate_0a,
  inp_0r, inp_0a, inp_0d,
  out_0r, out_0a, out_0d
);
  input activate_0r;
  output activate_0a;
  output inp_0r;
  input inp_0a;
  input [7:0] inp_0d;
  output out_0r;
  input out_0a;
  output [7:0] out_0d;
  assign activate_0a = out_0a;
  assign out_0r = inp_0a;
  assign inp_0r = activate_0r;
  assign out_0d[0] = inp_0d[0];
  assign out_0d[1] = inp_0d[1];
  assign out_0d[2] = inp_0d[2];
  assign out_0d[3] = inp_0d[3];
  assign out_0d[4] = inp_0d[4];
  assign out_0d[5] = inp_0d[5];
  assign out_0d[6] = inp_0d[6];
  assign out_0d[7] = inp_0d[7];
endmodule

module BrzFetch_16_s5_false (
  activate_0r, activate_0a,
  inp_0r, inp_0a, inp_0d,
  out_0r, out_0a, out_0d
);
  input activate_0r;
  output activate_0a;
  output inp_0r;
  input inp_0a;
  input [15:0] inp_0d;
  output out_0r;
  input out_0a;
  output [15:0] out_0d;
  assign activate_0a = out_0a;
  assign out_0r = inp_0a;
  assign inp_0r = activate_0r;
  assign out_0d[0] = inp_0d[0];
  assign out_0d[1] = inp_0d[1];
  assign out_0d[2] = inp_0d[2];
  assign out_0d[3] = inp_0d[3];
  assign out_0d[4] = inp_0d[4];
  assign out_0d[5] = inp_0d[5];
  assign out_0d[6] = inp_0d[6];
  assign out_0d[7] = inp_0d[7];
  assign out_0d[8] = inp_0d[8];
  assign out_0d[9] = inp_0d[9];
  assign out_0d[10] = inp_0d[10];
  assign out_0d[11] = inp_0d[11];
  assign out_0d[12] = inp_0d[12];
  assign out_0d[13] = inp_0d[13];
  assign out_0d[14] = inp_0d[14];
  assign out_0d[15] = inp_0d[15];
endmodule

module BrzFetch_17_s5_false (
  activate_0r, activate_0a,
  inp_0r, inp_0a, inp_0d,
  out_0r, out_0a, out_0d
);
  input activate_0r;
  output activate_0a;
  output inp_0r;
  input inp_0a;
  input [16:0] inp_0d;
  output out_0r;
  input out_0a;
  output [16:0] out_0d;
  assign activate_0a = out_0a;
  assign out_0r = inp_0a;
  assign inp_0r = activate_0r;
  assign out_0d[0] = inp_0d[0];
  assign out_0d[1] = inp_0d[1];
  assign out_0d[2] = inp_0d[2];
  assign out_0d[3] = inp_0d[3];
  assign out_0d[4] = inp_0d[4];
  assign out_0d[5] = inp_0d[5];
  assign out_0d[6] = inp_0d[6];
  assign out_0d[7] = inp_0d[7];
  assign out_0d[8] = inp_0d[8];
  assign out_0d[9] = inp_0d[9];
  assign out_0d[10] = inp_0d[10];
  assign out_0d[11] = inp_0d[11];
  assign out_0d[12] = inp_0d[12];
  assign out_0d[13] = inp_0d[13];
  assign out_0d[14] = inp_0d[14];
  assign out_0d[15] = inp_0d[15];
  assign out_0d[16] = inp_0d[16];
endmodule

module BrzLoop (
  activate_0r, activate_0a,
  activateOut_0r, activateOut_0a
);
  input activate_0r;
  output activate_0a;
  output activateOut_0r;
  input activateOut_0a;
  wire nReq_0n;
  wire gnd;
  GND gnd_cell_instance (gnd);
  IV I0 (nReq_0n, activate_0r);
  NR2 I1 (activateOut_0r, nReq_0n, activateOut_0a);
  assign activate_0a = gnd;
endmodule

module selem (
  Ar,
  Aa,
  Br,
  Ba
);
  input Ar;
  output Aa;
  output Br;
  input Ba;
  wire s_0n;
  NC2P I0 (s_0n, Ar, Ba);
  NR2 I1 (Aa, Ba, s_0n);
  AN2 I2 (Br, Ar, s_0n);
endmodule

module BrzSequence_2_s1_S (
  activate_0r, activate_0a,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a
);
  input activate_0r;
  output activate_0a;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  wire [1:0] sreq_0n;
  assign activate_0a = activateOut_1a;
  assign activateOut_1r = sreq_0n[1];
  assign sreq_0n[0] = activate_0r;
  selem I3 (sreq_0n[0], sreq_0n[1], activateOut_0r, activateOut_0a);
endmodule

module BrzSequence_19_s18_SSSSSSSSSSSSSSSSSS (
  activate_0r, activate_0a,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a,
  activateOut_2r, activateOut_2a,
  activateOut_3r, activateOut_3a,
  activateOut_4r, activateOut_4a,
  activateOut_5r, activateOut_5a,
  activateOut_6r, activateOut_6a,
  activateOut_7r, activateOut_7a,
  activateOut_8r, activateOut_8a,
  activateOut_9r, activateOut_9a,
  activateOut_10r, activateOut_10a,
  activateOut_11r, activateOut_11a,
  activateOut_12r, activateOut_12a,
  activateOut_13r, activateOut_13a,
  activateOut_14r, activateOut_14a,
  activateOut_15r, activateOut_15a,
  activateOut_16r, activateOut_16a,
  activateOut_17r, activateOut_17a,
  activateOut_18r, activateOut_18a
);
  input activate_0r;
  output activate_0a;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  output activateOut_2r;
  input activateOut_2a;
  output activateOut_3r;
  input activateOut_3a;
  output activateOut_4r;
  input activateOut_4a;
  output activateOut_5r;
  input activateOut_5a;
  output activateOut_6r;
  input activateOut_6a;
  output activateOut_7r;
  input activateOut_7a;
  output activateOut_8r;
  input activateOut_8a;
  output activateOut_9r;
  input activateOut_9a;
  output activateOut_10r;
  input activateOut_10a;
  output activateOut_11r;
  input activateOut_11a;
  output activateOut_12r;
  input activateOut_12a;
  output activateOut_13r;
  input activateOut_13a;
  output activateOut_14r;
  input activateOut_14a;
  output activateOut_15r;
  input activateOut_15a;
  output activateOut_16r;
  input activateOut_16a;
  output activateOut_17r;
  input activateOut_17a;
  output activateOut_18r;
  input activateOut_18a;
  wire [18:0] sreq_0n;
  assign activate_0a = activateOut_18a;
  assign activateOut_18r = sreq_0n[18];
  assign sreq_0n[0] = activate_0r;
  selem I3 (sreq_0n[17], sreq_0n[18], activateOut_17r, activateOut_17a);
  selem I4 (sreq_0n[16], sreq_0n[17], activateOut_16r, activateOut_16a);
  selem I5 (sreq_0n[15], sreq_0n[16], activateOut_15r, activateOut_15a);
  selem I6 (sreq_0n[14], sreq_0n[15], activateOut_14r, activateOut_14a);
  selem I7 (sreq_0n[13], sreq_0n[14], activateOut_13r, activateOut_13a);
  selem I8 (sreq_0n[12], sreq_0n[13], activateOut_12r, activateOut_12a);
  selem I9 (sreq_0n[11], sreq_0n[12], activateOut_11r, activateOut_11a);
  selem I10 (sreq_0n[10], sreq_0n[11], activateOut_10r, activateOut_10a);
  selem I11 (sreq_0n[9], sreq_0n[10], activateOut_9r, activateOut_9a);
  selem I12 (sreq_0n[8], sreq_0n[9], activateOut_8r, activateOut_8a);
  selem I13 (sreq_0n[7], sreq_0n[8], activateOut_7r, activateOut_7a);
  selem I14 (sreq_0n[6], sreq_0n[7], activateOut_6r, activateOut_6a);
  selem I15 (sreq_0n[5], sreq_0n[6], activateOut_5r, activateOut_5a);
  selem I16 (sreq_0n[4], sreq_0n[5], activateOut_4r, activateOut_4a);
  selem I17 (sreq_0n[3], sreq_0n[4], activateOut_3r, activateOut_3a);
  selem I18 (sreq_0n[2], sreq_0n[3], activateOut_2r, activateOut_2a);
  selem I19 (sreq_0n[1], sreq_0n[2], activateOut_1r, activateOut_1a);
  selem I20 (sreq_0n[0], sreq_0n[1], activateOut_0r, activateOut_0a);
endmodule

module BrzSlice_1_18_16 (
  out_0r, out_0a, out_0d,
  inp_0r, inp_0a, inp_0d
);
  input out_0r;
  output out_0a;
  output out_0d;
  output inp_0r;
  input inp_0a;
  input [17:0] inp_0d;
  assign inp_0r = out_0r;
  assign out_0a = inp_0a;
  assign out_0d = inp_0d[16];
endmodule

module BrzSlice_16_18_1 (
  out_0r, out_0a, out_0d,
  inp_0r, inp_0a, inp_0d
);
  input out_0r;
  output out_0a;
  output [15:0] out_0d;
  output inp_0r;
  input inp_0a;
  input [17:0] inp_0d;
  assign inp_0r = out_0r;
  assign out_0a = inp_0a;
  assign out_0d[0] = inp_0d[1];
  assign out_0d[1] = inp_0d[2];
  assign out_0d[2] = inp_0d[3];
  assign out_0d[3] = inp_0d[4];
  assign out_0d[4] = inp_0d[5];
  assign out_0d[5] = inp_0d[6];
  assign out_0d[6] = inp_0d[7];
  assign out_0d[7] = inp_0d[8];
  assign out_0d[8] = inp_0d[9];
  assign out_0d[9] = inp_0d[10];
  assign out_0d[10] = inp_0d[11];
  assign out_0d[11] = inp_0d[12];
  assign out_0d[12] = inp_0d[13];
  assign out_0d[13] = inp_0d[14];
  assign out_0d[14] = inp_0d[15];
  assign out_0d[15] = inp_0d[16];
endmodule

module BrzUnaryFunc_1_1_s6_Invert_s5_false (
  out_0r, out_0a, out_0d,
  inp_0r, inp_0a, inp_0d
);
  input out_0r;
  output out_0a;
  output out_0d;
  output inp_0r;
  input inp_0a;
  input inp_0d;
  wire nStart_0n;
  wire [1:0] nCv_0n;
  wire [1:0] c_0n;
  wire i_0n;
  wire j_0n;
  wire start_0n;
  wire done_0n;
  IV I0 (out_0d, inp_0d);
  assign done_0n = start_0n;
  assign out_0a = done_0n;
  assign start_0n = inp_0a;
  assign inp_0r = out_0r;
endmodule

module BrzUnaryFunc_8_8_s6_Negate_s4_true (
  out_0r, out_0a, out_0d,
  inp_0r, inp_0a, inp_0d
);
  input out_0r;
  output out_0a;
  output [7:0] out_0d;
  output inp_0r;
  input inp_0a;
  input [7:0] inp_0d;
  wire [1:0] internal_0n;
  wire nStart_0n;
  wire [8:0] nCv_0n;
  wire [8:0] c_0n;
  wire [7:0] i_0n;
  wire [7:0] j_0n;
  wire start_0n;
  wire done_0n;
  wire gnd;
  wire vcc;
  GND gnd_cell_instance (gnd);
  VCC vcc_cell_instance (vcc);
  NR4 I0 (internal_0n[0], nCv_0n[1], nCv_0n[2], nCv_0n[3], nCv_0n[4]);
  NR4 I1 (internal_0n[1], nCv_0n[5], nCv_0n[6], nCv_0n[7], nCv_0n[8]);
  AN2 I2 (done_0n, internal_0n[0], internal_0n[1]);
  balsa_fa I3 (nStart_0n, i_0n[0], j_0n[0], nCv_0n[0], c_0n[0], nCv_0n[1], c_0n[1], out_0d[0]);
  balsa_fa I4 (nStart_0n, i_0n[1], j_0n[1], nCv_0n[1], c_0n[1], nCv_0n[2], c_0n[2], out_0d[1]);
  balsa_fa I5 (nStart_0n, i_0n[2], j_0n[2], nCv_0n[2], c_0n[2], nCv_0n[3], c_0n[3], out_0d[2]);
  balsa_fa I6 (nStart_0n, i_0n[3], j_0n[3], nCv_0n[3], c_0n[3], nCv_0n[4], c_0n[4], out_0d[3]);
  balsa_fa I7 (nStart_0n, i_0n[4], j_0n[4], nCv_0n[4], c_0n[4], nCv_0n[5], c_0n[5], out_0d[4]);
  balsa_fa I8 (nStart_0n, i_0n[5], j_0n[5], nCv_0n[5], c_0n[5], nCv_0n[6], c_0n[6], out_0d[5]);
  balsa_fa I9 (nStart_0n, i_0n[6], j_0n[6], nCv_0n[6], c_0n[6], nCv_0n[7], c_0n[7], out_0d[6]);
  balsa_fa I10 (nStart_0n, i_0n[7], j_0n[7], nCv_0n[7], c_0n[7], nCv_0n[8], c_0n[8], out_0d[7]);
  assign c_0n[0] = vcc;
  assign j_0n[0] = gnd;
  assign j_0n[1] = gnd;
  assign j_0n[2] = gnd;
  assign j_0n[3] = gnd;
  assign j_0n[4] = gnd;
  assign j_0n[5] = gnd;
  assign j_0n[6] = gnd;
  assign j_0n[7] = gnd;
  assign nCv_0n[0] = nStart_0n;
  IV I21 (i_0n[0], inp_0d[0]);
  IV I22 (i_0n[1], inp_0d[1]);
  IV I23 (i_0n[2], inp_0d[2]);
  IV I24 (i_0n[3], inp_0d[3]);
  IV I25 (i_0n[4], inp_0d[4]);
  IV I26 (i_0n[5], inp_0d[5]);
  IV I27 (i_0n[6], inp_0d[6]);
  IV I28 (i_0n[7], inp_0d[7]);
  IV I29 (nStart_0n, start_0n);
  assign out_0a = done_0n;
  assign start_0n = inp_0a;
  assign inp_0r = out_0r;
endmodule

module BrzVariable_1_1_s0_ (
  write_0r, write_0a, write_0d,
  read_0r, read_0a, read_0d
);
  input write_0r;
  output write_0a;
  input write_0d;
  input read_0r;
  output read_0a;
  output read_0d;
  wire data_0n;
  wire nWriteReq_0n;
  wire bWriteReq_0n;
  wire nbWriteReq_0n;
  assign read_0a = read_0r;
  assign read_0d = data_0n;
  LD1 I2 (write_0d, bWriteReq_0n, data_0n);
  IV I3 (write_0a, nbWriteReq_0n);
  IV I4 (nbWriteReq_0n, bWriteReq_0n);
  IV I5 (bWriteReq_0n, nWriteReq_0n);
  IV I6 (nWriteReq_0n, write_0r);
endmodule

module BrzVariable_8_1_s0_ (
  write_0r, write_0a, write_0d,
  read_0r, read_0a, read_0d
);
  input write_0r;
  output write_0a;
  input [7:0] write_0d;
  input read_0r;
  output read_0a;
  output [7:0] read_0d;
  wire [7:0] data_0n;
  wire nWriteReq_0n;
  wire bWriteReq_0n;
  wire nbWriteReq_0n;
  assign read_0a = read_0r;
  assign read_0d[0] = data_0n[0];
  assign read_0d[1] = data_0n[1];
  assign read_0d[2] = data_0n[2];
  assign read_0d[3] = data_0n[3];
  assign read_0d[4] = data_0n[4];
  assign read_0d[5] = data_0n[5];
  assign read_0d[6] = data_0n[6];
  assign read_0d[7] = data_0n[7];
  LD1 I9 (write_0d[0], bWriteReq_0n, data_0n[0]);
  LD1 I10 (write_0d[1], bWriteReq_0n, data_0n[1]);
  LD1 I11 (write_0d[2], bWriteReq_0n, data_0n[2]);
  LD1 I12 (write_0d[3], bWriteReq_0n, data_0n[3]);
  LD1 I13 (write_0d[4], bWriteReq_0n, data_0n[4]);
  LD1 I14 (write_0d[5], bWriteReq_0n, data_0n[5]);
  LD1 I15 (write_0d[6], bWriteReq_0n, data_0n[6]);
  LD1 I16 (write_0d[7], bWriteReq_0n, data_0n[7]);
  IV I17 (write_0a, nbWriteReq_0n);
  IV I18 (nbWriteReq_0n, bWriteReq_0n);
  IV I19 (bWriteReq_0n, nWriteReq_0n);
  IV I20 (nWriteReq_0n, write_0r);
endmodule

module BrzVariable_8_2_s0_ (
  write_0r, write_0a, write_0d,
  read_0r, read_0a, read_0d,
  read_1r, read_1a, read_1d
);
  input write_0r;
  output write_0a;
  input [7:0] write_0d;
  input read_0r;
  output read_0a;
  output [7:0] read_0d;
  input read_1r;
  output read_1a;
  output [7:0] read_1d;
  wire [7:0] data_0n;
  wire nWriteReq_0n;
  wire bWriteReq_0n;
  wire nbWriteReq_0n;
  assign read_0a = read_0r;
  assign read_1a = read_1r;
  assign read_1d[0] = data_0n[0];
  assign read_1d[1] = data_0n[1];
  assign read_1d[2] = data_0n[2];
  assign read_1d[3] = data_0n[3];
  assign read_1d[4] = data_0n[4];
  assign read_1d[5] = data_0n[5];
  assign read_1d[6] = data_0n[6];
  assign read_1d[7] = data_0n[7];
  assign read_0d[0] = data_0n[0];
  assign read_0d[1] = data_0n[1];
  assign read_0d[2] = data_0n[2];
  assign read_0d[3] = data_0n[3];
  assign read_0d[4] = data_0n[4];
  assign read_0d[5] = data_0n[5];
  assign read_0d[6] = data_0n[6];
  assign read_0d[7] = data_0n[7];
  LD1 I18 (write_0d[0], bWriteReq_0n, data_0n[0]);
  LD1 I19 (write_0d[1], bWriteReq_0n, data_0n[1]);
  LD1 I20 (write_0d[2], bWriteReq_0n, data_0n[2]);
  LD1 I21 (write_0d[3], bWriteReq_0n, data_0n[3]);
  LD1 I22 (write_0d[4], bWriteReq_0n, data_0n[4]);
  LD1 I23 (write_0d[5], bWriteReq_0n, data_0n[5]);
  LD1 I24 (write_0d[6], bWriteReq_0n, data_0n[6]);
  LD1 I25 (write_0d[7], bWriteReq_0n, data_0n[7]);
  IV I26 (write_0a, nbWriteReq_0n);
  IV I27 (nbWriteReq_0n, bWriteReq_0n);
  IV I28 (bWriteReq_0n, nWriteReq_0n);
  IV I29 (nWriteReq_0n, write_0r);
endmodule

module BrzVariable_17_1_s0_ (
  write_0r, write_0a, write_0d,
  read_0r, read_0a, read_0d
);
  input write_0r;
  output write_0a;
  input [16:0] write_0d;
  input read_0r;
  output read_0a;
  output [16:0] read_0d;
  wire [16:0] data_0n;
  wire nWriteReq_0n;
  wire bWriteReq_0n;
  wire nbWriteReq_0n;
  assign read_0a = read_0r;
  assign read_0d[0] = data_0n[0];
  assign read_0d[1] = data_0n[1];
  assign read_0d[2] = data_0n[2];
  assign read_0d[3] = data_0n[3];
  assign read_0d[4] = data_0n[4];
  assign read_0d[5] = data_0n[5];
  assign read_0d[6] = data_0n[6];
  assign read_0d[7] = data_0n[7];
  assign read_0d[8] = data_0n[8];
  assign read_0d[9] = data_0n[9];
  assign read_0d[10] = data_0n[10];
  assign read_0d[11] = data_0n[11];
  assign read_0d[12] = data_0n[12];
  assign read_0d[13] = data_0n[13];
  assign read_0d[14] = data_0n[14];
  assign read_0d[15] = data_0n[15];
  assign read_0d[16] = data_0n[16];
  LD1 I18 (write_0d[0], bWriteReq_0n, data_0n[0]);
  LD1 I19 (write_0d[1], bWriteReq_0n, data_0n[1]);
  LD1 I20 (write_0d[2], bWriteReq_0n, data_0n[2]);
  LD1 I21 (write_0d[3], bWriteReq_0n, data_0n[3]);
  LD1 I22 (write_0d[4], bWriteReq_0n, data_0n[4]);
  LD1 I23 (write_0d[5], bWriteReq_0n, data_0n[5]);
  LD1 I24 (write_0d[6], bWriteReq_0n, data_0n[6]);
  LD1 I25 (write_0d[7], bWriteReq_0n, data_0n[7]);
  LD1 I26 (write_0d[8], bWriteReq_0n, data_0n[8]);
  LD1 I27 (write_0d[9], bWriteReq_0n, data_0n[9]);
  LD1 I28 (write_0d[10], bWriteReq_0n, data_0n[10]);
  LD1 I29 (write_0d[11], bWriteReq_0n, data_0n[11]);
  LD1 I30 (write_0d[12], bWriteReq_0n, data_0n[12]);
  LD1 I31 (write_0d[13], bWriteReq_0n, data_0n[13]);
  LD1 I32 (write_0d[14], bWriteReq_0n, data_0n[14]);
  LD1 I33 (write_0d[15], bWriteReq_0n, data_0n[15]);
  LD1 I34 (write_0d[16], bWriteReq_0n, data_0n[16]);
  IV I35 (write_0a, nbWriteReq_0n);
  IV I36 (nbWriteReq_0n, bWriteReq_0n);
  IV I37 (bWriteReq_0n, nWriteReq_0n);
  IV I38 (nWriteReq_0n, write_0r);
endmodule

module BrzVariable_17_16_s0_ (
  write_0r, write_0a, write_0d,
  read_0r, read_0a, read_0d,
  read_1r, read_1a, read_1d,
  read_2r, read_2a, read_2d,
  read_3r, read_3a, read_3d,
  read_4r, read_4a, read_4d,
  read_5r, read_5a, read_5d,
  read_6r, read_6a, read_6d,
  read_7r, read_7a, read_7d,
  read_8r, read_8a, read_8d,
  read_9r, read_9a, read_9d,
  read_10r, read_10a, read_10d,
  read_11r, read_11a, read_11d,
  read_12r, read_12a, read_12d,
  read_13r, read_13a, read_13d,
  read_14r, read_14a, read_14d,
  read_15r, read_15a, read_15d
);
  input write_0r;
  output write_0a;
  input [16:0] write_0d;
  input read_0r;
  output read_0a;
  output [16:0] read_0d;
  input read_1r;
  output read_1a;
  output [16:0] read_1d;
  input read_2r;
  output read_2a;
  output [16:0] read_2d;
  input read_3r;
  output read_3a;
  output [16:0] read_3d;
  input read_4r;
  output read_4a;
  output [16:0] read_4d;
  input read_5r;
  output read_5a;
  output [16:0] read_5d;
  input read_6r;
  output read_6a;
  output [16:0] read_6d;
  input read_7r;
  output read_7a;
  output [16:0] read_7d;
  input read_8r;
  output read_8a;
  output [16:0] read_8d;
  input read_9r;
  output read_9a;
  output [16:0] read_9d;
  input read_10r;
  output read_10a;
  output [16:0] read_10d;
  input read_11r;
  output read_11a;
  output [16:0] read_11d;
  input read_12r;
  output read_12a;
  output [16:0] read_12d;
  input read_13r;
  output read_13a;
  output [16:0] read_13d;
  input read_14r;
  output read_14a;
  output [16:0] read_14d;
  input read_15r;
  output read_15a;
  output [16:0] read_15d;
  wire [16:0] data_0n;
  wire nWriteReq_0n;
  wire bWriteReq_0n;
  wire nbWriteReq_0n;
  assign read_0a = read_0r;
  assign read_1a = read_1r;
  assign read_2a = read_2r;
  assign read_3a = read_3r;
  assign read_4a = read_4r;
  assign read_5a = read_5r;
  assign read_6a = read_6r;
  assign read_7a = read_7r;
  assign read_8a = read_8r;
  assign read_9a = read_9r;
  assign read_10a = read_10r;
  assign read_11a = read_11r;
  assign read_12a = read_12r;
  assign read_13a = read_13r;
  assign read_14a = read_14r;
  assign read_15a = read_15r;
  assign read_15d[0] = data_0n[0];
  assign read_15d[1] = data_0n[1];
  assign read_15d[2] = data_0n[2];
  assign read_15d[3] = data_0n[3];
  assign read_15d[4] = data_0n[4];
  assign read_15d[5] = data_0n[5];
  assign read_15d[6] = data_0n[6];
  assign read_15d[7] = data_0n[7];
  assign read_15d[8] = data_0n[8];
  assign read_15d[9] = data_0n[9];
  assign read_15d[10] = data_0n[10];
  assign read_15d[11] = data_0n[11];
  assign read_15d[12] = data_0n[12];
  assign read_15d[13] = data_0n[13];
  assign read_15d[14] = data_0n[14];
  assign read_15d[15] = data_0n[15];
  assign read_15d[16] = data_0n[16];
  assign read_14d[0] = data_0n[0];
  assign read_14d[1] = data_0n[1];
  assign read_14d[2] = data_0n[2];
  assign read_14d[3] = data_0n[3];
  assign read_14d[4] = data_0n[4];
  assign read_14d[5] = data_0n[5];
  assign read_14d[6] = data_0n[6];
  assign read_14d[7] = data_0n[7];
  assign read_14d[8] = data_0n[8];
  assign read_14d[9] = data_0n[9];
  assign read_14d[10] = data_0n[10];
  assign read_14d[11] = data_0n[11];
  assign read_14d[12] = data_0n[12];
  assign read_14d[13] = data_0n[13];
  assign read_14d[14] = data_0n[14];
  assign read_14d[15] = data_0n[15];
  assign read_14d[16] = data_0n[16];
  assign read_13d[0] = data_0n[0];
  assign read_13d[1] = data_0n[1];
  assign read_13d[2] = data_0n[2];
  assign read_13d[3] = data_0n[3];
  assign read_13d[4] = data_0n[4];
  assign read_13d[5] = data_0n[5];
  assign read_13d[6] = data_0n[6];
  assign read_13d[7] = data_0n[7];
  assign read_13d[8] = data_0n[8];
  assign read_13d[9] = data_0n[9];
  assign read_13d[10] = data_0n[10];
  assign read_13d[11] = data_0n[11];
  assign read_13d[12] = data_0n[12];
  assign read_13d[13] = data_0n[13];
  assign read_13d[14] = data_0n[14];
  assign read_13d[15] = data_0n[15];
  assign read_13d[16] = data_0n[16];
  assign read_12d[0] = data_0n[0];
  assign read_12d[1] = data_0n[1];
  assign read_12d[2] = data_0n[2];
  assign read_12d[3] = data_0n[3];
  assign read_12d[4] = data_0n[4];
  assign read_12d[5] = data_0n[5];
  assign read_12d[6] = data_0n[6];
  assign read_12d[7] = data_0n[7];
  assign read_12d[8] = data_0n[8];
  assign read_12d[9] = data_0n[9];
  assign read_12d[10] = data_0n[10];
  assign read_12d[11] = data_0n[11];
  assign read_12d[12] = data_0n[12];
  assign read_12d[13] = data_0n[13];
  assign read_12d[14] = data_0n[14];
  assign read_12d[15] = data_0n[15];
  assign read_12d[16] = data_0n[16];
  assign read_11d[0] = data_0n[0];
  assign read_11d[1] = data_0n[1];
  assign read_11d[2] = data_0n[2];
  assign read_11d[3] = data_0n[3];
  assign read_11d[4] = data_0n[4];
  assign read_11d[5] = data_0n[5];
  assign read_11d[6] = data_0n[6];
  assign read_11d[7] = data_0n[7];
  assign read_11d[8] = data_0n[8];
  assign read_11d[9] = data_0n[9];
  assign read_11d[10] = data_0n[10];
  assign read_11d[11] = data_0n[11];
  assign read_11d[12] = data_0n[12];
  assign read_11d[13] = data_0n[13];
  assign read_11d[14] = data_0n[14];
  assign read_11d[15] = data_0n[15];
  assign read_11d[16] = data_0n[16];
  assign read_10d[0] = data_0n[0];
  assign read_10d[1] = data_0n[1];
  assign read_10d[2] = data_0n[2];
  assign read_10d[3] = data_0n[3];
  assign read_10d[4] = data_0n[4];
  assign read_10d[5] = data_0n[5];
  assign read_10d[6] = data_0n[6];
  assign read_10d[7] = data_0n[7];
  assign read_10d[8] = data_0n[8];
  assign read_10d[9] = data_0n[9];
  assign read_10d[10] = data_0n[10];
  assign read_10d[11] = data_0n[11];
  assign read_10d[12] = data_0n[12];
  assign read_10d[13] = data_0n[13];
  assign read_10d[14] = data_0n[14];
  assign read_10d[15] = data_0n[15];
  assign read_10d[16] = data_0n[16];
  assign read_9d[0] = data_0n[0];
  assign read_9d[1] = data_0n[1];
  assign read_9d[2] = data_0n[2];
  assign read_9d[3] = data_0n[3];
  assign read_9d[4] = data_0n[4];
  assign read_9d[5] = data_0n[5];
  assign read_9d[6] = data_0n[6];
  assign read_9d[7] = data_0n[7];
  assign read_9d[8] = data_0n[8];
  assign read_9d[9] = data_0n[9];
  assign read_9d[10] = data_0n[10];
  assign read_9d[11] = data_0n[11];
  assign read_9d[12] = data_0n[12];
  assign read_9d[13] = data_0n[13];
  assign read_9d[14] = data_0n[14];
  assign read_9d[15] = data_0n[15];
  assign read_9d[16] = data_0n[16];
  assign read_8d[0] = data_0n[0];
  assign read_8d[1] = data_0n[1];
  assign read_8d[2] = data_0n[2];
  assign read_8d[3] = data_0n[3];
  assign read_8d[4] = data_0n[4];
  assign read_8d[5] = data_0n[5];
  assign read_8d[6] = data_0n[6];
  assign read_8d[7] = data_0n[7];
  assign read_8d[8] = data_0n[8];
  assign read_8d[9] = data_0n[9];
  assign read_8d[10] = data_0n[10];
  assign read_8d[11] = data_0n[11];
  assign read_8d[12] = data_0n[12];
  assign read_8d[13] = data_0n[13];
  assign read_8d[14] = data_0n[14];
  assign read_8d[15] = data_0n[15];
  assign read_8d[16] = data_0n[16];
  assign read_7d[0] = data_0n[0];
  assign read_7d[1] = data_0n[1];
  assign read_7d[2] = data_0n[2];
  assign read_7d[3] = data_0n[3];
  assign read_7d[4] = data_0n[4];
  assign read_7d[5] = data_0n[5];
  assign read_7d[6] = data_0n[6];
  assign read_7d[7] = data_0n[7];
  assign read_7d[8] = data_0n[8];
  assign read_7d[9] = data_0n[9];
  assign read_7d[10] = data_0n[10];
  assign read_7d[11] = data_0n[11];
  assign read_7d[12] = data_0n[12];
  assign read_7d[13] = data_0n[13];
  assign read_7d[14] = data_0n[14];
  assign read_7d[15] = data_0n[15];
  assign read_7d[16] = data_0n[16];
  assign read_6d[0] = data_0n[0];
  assign read_6d[1] = data_0n[1];
  assign read_6d[2] = data_0n[2];
  assign read_6d[3] = data_0n[3];
  assign read_6d[4] = data_0n[4];
  assign read_6d[5] = data_0n[5];
  assign read_6d[6] = data_0n[6];
  assign read_6d[7] = data_0n[7];
  assign read_6d[8] = data_0n[8];
  assign read_6d[9] = data_0n[9];
  assign read_6d[10] = data_0n[10];
  assign read_6d[11] = data_0n[11];
  assign read_6d[12] = data_0n[12];
  assign read_6d[13] = data_0n[13];
  assign read_6d[14] = data_0n[14];
  assign read_6d[15] = data_0n[15];
  assign read_6d[16] = data_0n[16];
  assign read_5d[0] = data_0n[0];
  assign read_5d[1] = data_0n[1];
  assign read_5d[2] = data_0n[2];
  assign read_5d[3] = data_0n[3];
  assign read_5d[4] = data_0n[4];
  assign read_5d[5] = data_0n[5];
  assign read_5d[6] = data_0n[6];
  assign read_5d[7] = data_0n[7];
  assign read_5d[8] = data_0n[8];
  assign read_5d[9] = data_0n[9];
  assign read_5d[10] = data_0n[10];
  assign read_5d[11] = data_0n[11];
  assign read_5d[12] = data_0n[12];
  assign read_5d[13] = data_0n[13];
  assign read_5d[14] = data_0n[14];
  assign read_5d[15] = data_0n[15];
  assign read_5d[16] = data_0n[16];
  assign read_4d[0] = data_0n[0];
  assign read_4d[1] = data_0n[1];
  assign read_4d[2] = data_0n[2];
  assign read_4d[3] = data_0n[3];
  assign read_4d[4] = data_0n[4];
  assign read_4d[5] = data_0n[5];
  assign read_4d[6] = data_0n[6];
  assign read_4d[7] = data_0n[7];
  assign read_4d[8] = data_0n[8];
  assign read_4d[9] = data_0n[9];
  assign read_4d[10] = data_0n[10];
  assign read_4d[11] = data_0n[11];
  assign read_4d[12] = data_0n[12];
  assign read_4d[13] = data_0n[13];
  assign read_4d[14] = data_0n[14];
  assign read_4d[15] = data_0n[15];
  assign read_4d[16] = data_0n[16];
  assign read_3d[0] = data_0n[0];
  assign read_3d[1] = data_0n[1];
  assign read_3d[2] = data_0n[2];
  assign read_3d[3] = data_0n[3];
  assign read_3d[4] = data_0n[4];
  assign read_3d[5] = data_0n[5];
  assign read_3d[6] = data_0n[6];
  assign read_3d[7] = data_0n[7];
  assign read_3d[8] = data_0n[8];
  assign read_3d[9] = data_0n[9];
  assign read_3d[10] = data_0n[10];
  assign read_3d[11] = data_0n[11];
  assign read_3d[12] = data_0n[12];
  assign read_3d[13] = data_0n[13];
  assign read_3d[14] = data_0n[14];
  assign read_3d[15] = data_0n[15];
  assign read_3d[16] = data_0n[16];
  assign read_2d[0] = data_0n[0];
  assign read_2d[1] = data_0n[1];
  assign read_2d[2] = data_0n[2];
  assign read_2d[3] = data_0n[3];
  assign read_2d[4] = data_0n[4];
  assign read_2d[5] = data_0n[5];
  assign read_2d[6] = data_0n[6];
  assign read_2d[7] = data_0n[7];
  assign read_2d[8] = data_0n[8];
  assign read_2d[9] = data_0n[9];
  assign read_2d[10] = data_0n[10];
  assign read_2d[11] = data_0n[11];
  assign read_2d[12] = data_0n[12];
  assign read_2d[13] = data_0n[13];
  assign read_2d[14] = data_0n[14];
  assign read_2d[15] = data_0n[15];
  assign read_2d[16] = data_0n[16];
  assign read_1d[0] = data_0n[0];
  assign read_1d[1] = data_0n[1];
  assign read_1d[2] = data_0n[2];
  assign read_1d[3] = data_0n[3];
  assign read_1d[4] = data_0n[4];
  assign read_1d[5] = data_0n[5];
  assign read_1d[6] = data_0n[6];
  assign read_1d[7] = data_0n[7];
  assign read_1d[8] = data_0n[8];
  assign read_1d[9] = data_0n[9];
  assign read_1d[10] = data_0n[10];
  assign read_1d[11] = data_0n[11];
  assign read_1d[12] = data_0n[12];
  assign read_1d[13] = data_0n[13];
  assign read_1d[14] = data_0n[14];
  assign read_1d[15] = data_0n[15];
  assign read_1d[16] = data_0n[16];
  assign read_0d[0] = data_0n[0];
  assign read_0d[1] = data_0n[1];
  assign read_0d[2] = data_0n[2];
  assign read_0d[3] = data_0n[3];
  assign read_0d[4] = data_0n[4];
  assign read_0d[5] = data_0n[5];
  assign read_0d[6] = data_0n[6];
  assign read_0d[7] = data_0n[7];
  assign read_0d[8] = data_0n[8];
  assign read_0d[9] = data_0n[9];
  assign read_0d[10] = data_0n[10];
  assign read_0d[11] = data_0n[11];
  assign read_0d[12] = data_0n[12];
  assign read_0d[13] = data_0n[13];
  assign read_0d[14] = data_0n[14];
  assign read_0d[15] = data_0n[15];
  assign read_0d[16] = data_0n[16];
  LD1 I288 (write_0d[0], bWriteReq_0n, data_0n[0]);
  LD1 I289 (write_0d[1], bWriteReq_0n, data_0n[1]);
  LD1 I290 (write_0d[2], bWriteReq_0n, data_0n[2]);
  LD1 I291 (write_0d[3], bWriteReq_0n, data_0n[3]);
  LD1 I292 (write_0d[4], bWriteReq_0n, data_0n[4]);
  LD1 I293 (write_0d[5], bWriteReq_0n, data_0n[5]);
  LD1 I294 (write_0d[6], bWriteReq_0n, data_0n[6]);
  LD1 I295 (write_0d[7], bWriteReq_0n, data_0n[7]);
  LD1 I296 (write_0d[8], bWriteReq_0n, data_0n[8]);
  LD1 I297 (write_0d[9], bWriteReq_0n, data_0n[9]);
  LD1 I298 (write_0d[10], bWriteReq_0n, data_0n[10]);
  LD1 I299 (write_0d[11], bWriteReq_0n, data_0n[11]);
  LD1 I300 (write_0d[12], bWriteReq_0n, data_0n[12]);
  LD1 I301 (write_0d[13], bWriteReq_0n, data_0n[13]);
  LD1 I302 (write_0d[14], bWriteReq_0n, data_0n[14]);
  LD1 I303 (write_0d[15], bWriteReq_0n, data_0n[15]);
  LD1 I304 (write_0d[16], bWriteReq_0n, data_0n[16]);
  IV I305 (write_0a, nbWriteReq_0n);
  IV I306 (nbWriteReq_0n, bWriteReq_0n);
  IV I307 (bWriteReq_0n, nWriteReq_0n);
  IV I308 (nWriteReq_0n, write_0r);
endmodule

module BrzVariable_17_81_s657_1_2e_2e1_3b0_2e_2e0_m6m (
  write_0r, write_0a, write_0d,
  read_0r, read_0a, read_0d,
  read_1r, read_1a, read_1d,
  read_2r, read_2a, read_2d,
  read_3r, read_3a, read_3d,
  read_4r, read_4a, read_4d,
  read_5r, read_5a, read_5d,
  read_6r, read_6a, read_6d,
  read_7r, read_7a, read_7d,
  read_8r, read_8a, read_8d,
  read_9r, read_9a, read_9d,
  read_10r, read_10a, read_10d,
  read_11r, read_11a, read_11d,
  read_12r, read_12a, read_12d,
  read_13r, read_13a, read_13d,
  read_14r, read_14a, read_14d,
  read_15r, read_15a, read_15d,
  read_16r, read_16a, read_16d,
  read_17r, read_17a, read_17d,
  read_18r, read_18a, read_18d,
  read_19r, read_19a, read_19d,
  read_20r, read_20a, read_20d,
  read_21r, read_21a, read_21d,
  read_22r, read_22a, read_22d,
  read_23r, read_23a, read_23d,
  read_24r, read_24a, read_24d,
  read_25r, read_25a, read_25d,
  read_26r, read_26a, read_26d,
  read_27r, read_27a, read_27d,
  read_28r, read_28a, read_28d,
  read_29r, read_29a, read_29d,
  read_30r, read_30a, read_30d,
  read_31r, read_31a, read_31d,
  read_32r, read_32a, read_32d,
  read_33r, read_33a, read_33d,
  read_34r, read_34a, read_34d,
  read_35r, read_35a, read_35d,
  read_36r, read_36a, read_36d,
  read_37r, read_37a, read_37d,
  read_38r, read_38a, read_38d,
  read_39r, read_39a, read_39d,
  read_40r, read_40a, read_40d,
  read_41r, read_41a, read_41d,
  read_42r, read_42a, read_42d,
  read_43r, read_43a, read_43d,
  read_44r, read_44a, read_44d,
  read_45r, read_45a, read_45d,
  read_46r, read_46a, read_46d,
  read_47r, read_47a, read_47d,
  read_48r, read_48a, read_48d,
  read_49r, read_49a, read_49d,
  read_50r, read_50a, read_50d,
  read_51r, read_51a, read_51d,
  read_52r, read_52a, read_52d,
  read_53r, read_53a, read_53d,
  read_54r, read_54a, read_54d,
  read_55r, read_55a, read_55d,
  read_56r, read_56a, read_56d,
  read_57r, read_57a, read_57d,
  read_58r, read_58a, read_58d,
  read_59r, read_59a, read_59d,
  read_60r, read_60a, read_60d,
  read_61r, read_61a, read_61d,
  read_62r, read_62a, read_62d,
  read_63r, read_63a, read_63d,
  read_64r, read_64a, read_64d,
  read_65r, read_65a, read_65d,
  read_66r, read_66a, read_66d,
  read_67r, read_67a, read_67d,
  read_68r, read_68a, read_68d,
  read_69r, read_69a, read_69d,
  read_70r, read_70a, read_70d,
  read_71r, read_71a, read_71d,
  read_72r, read_72a, read_72d,
  read_73r, read_73a, read_73d,
  read_74r, read_74a, read_74d,
  read_75r, read_75a, read_75d,
  read_76r, read_76a, read_76d,
  read_77r, read_77a, read_77d,
  read_78r, read_78a, read_78d,
  read_79r, read_79a, read_79d,
  read_80r, read_80a, read_80d
);
  input write_0r;
  output write_0a;
  input [16:0] write_0d;
  input read_0r;
  output read_0a;
  output read_0d;
  input read_1r;
  output read_1a;
  output read_1d;
  input read_2r;
  output read_2a;
  output read_2d;
  input read_3r;
  output read_3a;
  output read_3d;
  input read_4r;
  output read_4a;
  output [16:0] read_4d;
  input read_5r;
  output read_5a;
  output [16:0] read_5d;
  input read_6r;
  output read_6a;
  output [16:0] read_6d;
  input read_7r;
  output read_7a;
  output [16:0] read_7d;
  input read_8r;
  output read_8a;
  output [15:0] read_8d;
  input read_9r;
  output read_9a;
  output read_9d;
  input read_10r;
  output read_10a;
  output read_10d;
  input read_11r;
  output read_11a;
  output read_11d;
  input read_12r;
  output read_12a;
  output read_12d;
  input read_13r;
  output read_13a;
  output read_13d;
  input read_14r;
  output read_14a;
  output [16:0] read_14d;
  input read_15r;
  output read_15a;
  output [16:0] read_15d;
  input read_16r;
  output read_16a;
  output [16:0] read_16d;
  input read_17r;
  output read_17a;
  output [16:0] read_17d;
  input read_18r;
  output read_18a;
  output [15:0] read_18d;
  input read_19r;
  output read_19a;
  output read_19d;
  input read_20r;
  output read_20a;
  output read_20d;
  input read_21r;
  output read_21a;
  output read_21d;
  input read_22r;
  output read_22a;
  output read_22d;
  input read_23r;
  output read_23a;
  output read_23d;
  input read_24r;
  output read_24a;
  output [16:0] read_24d;
  input read_25r;
  output read_25a;
  output [16:0] read_25d;
  input read_26r;
  output read_26a;
  output [16:0] read_26d;
  input read_27r;
  output read_27a;
  output [16:0] read_27d;
  input read_28r;
  output read_28a;
  output [15:0] read_28d;
  input read_29r;
  output read_29a;
  output read_29d;
  input read_30r;
  output read_30a;
  output read_30d;
  input read_31r;
  output read_31a;
  output read_31d;
  input read_32r;
  output read_32a;
  output read_32d;
  input read_33r;
  output read_33a;
  output read_33d;
  input read_34r;
  output read_34a;
  output [16:0] read_34d;
  input read_35r;
  output read_35a;
  output [16:0] read_35d;
  input read_36r;
  output read_36a;
  output [16:0] read_36d;
  input read_37r;
  output read_37a;
  output [16:0] read_37d;
  input read_38r;
  output read_38a;
  output [15:0] read_38d;
  input read_39r;
  output read_39a;
  output read_39d;
  input read_40r;
  output read_40a;
  output read_40d;
  input read_41r;
  output read_41a;
  output read_41d;
  input read_42r;
  output read_42a;
  output read_42d;
  input read_43r;
  output read_43a;
  output read_43d;
  input read_44r;
  output read_44a;
  output [16:0] read_44d;
  input read_45r;
  output read_45a;
  output [16:0] read_45d;
  input read_46r;
  output read_46a;
  output [16:0] read_46d;
  input read_47r;
  output read_47a;
  output [16:0] read_47d;
  input read_48r;
  output read_48a;
  output [15:0] read_48d;
  input read_49r;
  output read_49a;
  output read_49d;
  input read_50r;
  output read_50a;
  output read_50d;
  input read_51r;
  output read_51a;
  output read_51d;
  input read_52r;
  output read_52a;
  output read_52d;
  input read_53r;
  output read_53a;
  output read_53d;
  input read_54r;
  output read_54a;
  output [16:0] read_54d;
  input read_55r;
  output read_55a;
  output [16:0] read_55d;
  input read_56r;
  output read_56a;
  output [16:0] read_56d;
  input read_57r;
  output read_57a;
  output [16:0] read_57d;
  input read_58r;
  output read_58a;
  output [15:0] read_58d;
  input read_59r;
  output read_59a;
  output read_59d;
  input read_60r;
  output read_60a;
  output read_60d;
  input read_61r;
  output read_61a;
  output read_61d;
  input read_62r;
  output read_62a;
  output read_62d;
  input read_63r;
  output read_63a;
  output read_63d;
  input read_64r;
  output read_64a;
  output [16:0] read_64d;
  input read_65r;
  output read_65a;
  output [16:0] read_65d;
  input read_66r;
  output read_66a;
  output [16:0] read_66d;
  input read_67r;
  output read_67a;
  output [16:0] read_67d;
  input read_68r;
  output read_68a;
  output [15:0] read_68d;
  input read_69r;
  output read_69a;
  output read_69d;
  input read_70r;
  output read_70a;
  output read_70d;
  input read_71r;
  output read_71a;
  output read_71d;
  input read_72r;
  output read_72a;
  output read_72d;
  input read_73r;
  output read_73a;
  output read_73d;
  input read_74r;
  output read_74a;
  output [16:0] read_74d;
  input read_75r;
  output read_75a;
  output [16:0] read_75d;
  input read_76r;
  output read_76a;
  output [16:0] read_76d;
  input read_77r;
  output read_77a;
  output [16:0] read_77d;
  input read_78r;
  output read_78a;
  output [15:0] read_78d;
  input read_79r;
  output read_79a;
  output read_79d;
  input read_80r;
  output read_80a;
  output [15:0] read_80d;
  wire [16:0] data_0n;
  wire nWriteReq_0n;
  wire bWriteReq_0n;
  wire nbWriteReq_0n;
  assign read_0a = read_0r;
  assign read_1a = read_1r;
  assign read_2a = read_2r;
  assign read_3a = read_3r;
  assign read_4a = read_4r;
  assign read_5a = read_5r;
  assign read_6a = read_6r;
  assign read_7a = read_7r;
  assign read_8a = read_8r;
  assign read_9a = read_9r;
  assign read_10a = read_10r;
  assign read_11a = read_11r;
  assign read_12a = read_12r;
  assign read_13a = read_13r;
  assign read_14a = read_14r;
  assign read_15a = read_15r;
  assign read_16a = read_16r;
  assign read_17a = read_17r;
  assign read_18a = read_18r;
  assign read_19a = read_19r;
  assign read_20a = read_20r;
  assign read_21a = read_21r;
  assign read_22a = read_22r;
  assign read_23a = read_23r;
  assign read_24a = read_24r;
  assign read_25a = read_25r;
  assign read_26a = read_26r;
  assign read_27a = read_27r;
  assign read_28a = read_28r;
  assign read_29a = read_29r;
  assign read_30a = read_30r;
  assign read_31a = read_31r;
  assign read_32a = read_32r;
  assign read_33a = read_33r;
  assign read_34a = read_34r;
  assign read_35a = read_35r;
  assign read_36a = read_36r;
  assign read_37a = read_37r;
  assign read_38a = read_38r;
  assign read_39a = read_39r;
  assign read_40a = read_40r;
  assign read_41a = read_41r;
  assign read_42a = read_42r;
  assign read_43a = read_43r;
  assign read_44a = read_44r;
  assign read_45a = read_45r;
  assign read_46a = read_46r;
  assign read_47a = read_47r;
  assign read_48a = read_48r;
  assign read_49a = read_49r;
  assign read_50a = read_50r;
  assign read_51a = read_51r;
  assign read_52a = read_52r;
  assign read_53a = read_53r;
  assign read_54a = read_54r;
  assign read_55a = read_55r;
  assign read_56a = read_56r;
  assign read_57a = read_57r;
  assign read_58a = read_58r;
  assign read_59a = read_59r;
  assign read_60a = read_60r;
  assign read_61a = read_61r;
  assign read_62a = read_62r;
  assign read_63a = read_63r;
  assign read_64a = read_64r;
  assign read_65a = read_65r;
  assign read_66a = read_66r;
  assign read_67a = read_67r;
  assign read_68a = read_68r;
  assign read_69a = read_69r;
  assign read_70a = read_70r;
  assign read_71a = read_71r;
  assign read_72a = read_72r;
  assign read_73a = read_73r;
  assign read_74a = read_74r;
  assign read_75a = read_75r;
  assign read_76a = read_76r;
  assign read_77a = read_77r;
  assign read_78a = read_78r;
  assign read_79a = read_79r;
  assign read_80a = read_80r;
  assign read_80d[0] = data_0n[1];
  assign read_80d[1] = data_0n[2];
  assign read_80d[2] = data_0n[3];
  assign read_80d[3] = data_0n[4];
  assign read_80d[4] = data_0n[5];
  assign read_80d[5] = data_0n[6];
  assign read_80d[6] = data_0n[7];
  assign read_80d[7] = data_0n[8];
  assign read_80d[8] = data_0n[9];
  assign read_80d[9] = data_0n[10];
  assign read_80d[10] = data_0n[11];
  assign read_80d[11] = data_0n[12];
  assign read_80d[12] = data_0n[13];
  assign read_80d[13] = data_0n[14];
  assign read_80d[14] = data_0n[15];
  assign read_80d[15] = data_0n[16];
  assign read_79d = data_0n[16];
  assign read_78d[0] = data_0n[1];
  assign read_78d[1] = data_0n[2];
  assign read_78d[2] = data_0n[3];
  assign read_78d[3] = data_0n[4];
  assign read_78d[4] = data_0n[5];
  assign read_78d[5] = data_0n[6];
  assign read_78d[6] = data_0n[7];
  assign read_78d[7] = data_0n[8];
  assign read_78d[8] = data_0n[9];
  assign read_78d[9] = data_0n[10];
  assign read_78d[10] = data_0n[11];
  assign read_78d[11] = data_0n[12];
  assign read_78d[12] = data_0n[13];
  assign read_78d[13] = data_0n[14];
  assign read_78d[14] = data_0n[15];
  assign read_78d[15] = data_0n[16];
  assign read_77d[0] = data_0n[0];
  assign read_77d[1] = data_0n[1];
  assign read_77d[2] = data_0n[2];
  assign read_77d[3] = data_0n[3];
  assign read_77d[4] = data_0n[4];
  assign read_77d[5] = data_0n[5];
  assign read_77d[6] = data_0n[6];
  assign read_77d[7] = data_0n[7];
  assign read_77d[8] = data_0n[8];
  assign read_77d[9] = data_0n[9];
  assign read_77d[10] = data_0n[10];
  assign read_77d[11] = data_0n[11];
  assign read_77d[12] = data_0n[12];
  assign read_77d[13] = data_0n[13];
  assign read_77d[14] = data_0n[14];
  assign read_77d[15] = data_0n[15];
  assign read_77d[16] = data_0n[16];
  assign read_76d[0] = data_0n[0];
  assign read_76d[1] = data_0n[1];
  assign read_76d[2] = data_0n[2];
  assign read_76d[3] = data_0n[3];
  assign read_76d[4] = data_0n[4];
  assign read_76d[5] = data_0n[5];
  assign read_76d[6] = data_0n[6];
  assign read_76d[7] = data_0n[7];
  assign read_76d[8] = data_0n[8];
  assign read_76d[9] = data_0n[9];
  assign read_76d[10] = data_0n[10];
  assign read_76d[11] = data_0n[11];
  assign read_76d[12] = data_0n[12];
  assign read_76d[13] = data_0n[13];
  assign read_76d[14] = data_0n[14];
  assign read_76d[15] = data_0n[15];
  assign read_76d[16] = data_0n[16];
  assign read_75d[0] = data_0n[0];
  assign read_75d[1] = data_0n[1];
  assign read_75d[2] = data_0n[2];
  assign read_75d[3] = data_0n[3];
  assign read_75d[4] = data_0n[4];
  assign read_75d[5] = data_0n[5];
  assign read_75d[6] = data_0n[6];
  assign read_75d[7] = data_0n[7];
  assign read_75d[8] = data_0n[8];
  assign read_75d[9] = data_0n[9];
  assign read_75d[10] = data_0n[10];
  assign read_75d[11] = data_0n[11];
  assign read_75d[12] = data_0n[12];
  assign read_75d[13] = data_0n[13];
  assign read_75d[14] = data_0n[14];
  assign read_75d[15] = data_0n[15];
  assign read_75d[16] = data_0n[16];
  assign read_74d[0] = data_0n[0];
  assign read_74d[1] = data_0n[1];
  assign read_74d[2] = data_0n[2];
  assign read_74d[3] = data_0n[3];
  assign read_74d[4] = data_0n[4];
  assign read_74d[5] = data_0n[5];
  assign read_74d[6] = data_0n[6];
  assign read_74d[7] = data_0n[7];
  assign read_74d[8] = data_0n[8];
  assign read_74d[9] = data_0n[9];
  assign read_74d[10] = data_0n[10];
  assign read_74d[11] = data_0n[11];
  assign read_74d[12] = data_0n[12];
  assign read_74d[13] = data_0n[13];
  assign read_74d[14] = data_0n[14];
  assign read_74d[15] = data_0n[15];
  assign read_74d[16] = data_0n[16];
  assign read_73d = data_0n[0];
  assign read_72d = data_0n[1];
  assign read_71d = data_0n[0];
  assign read_70d = data_0n[1];
  assign read_69d = data_0n[16];
  assign read_68d[0] = data_0n[1];
  assign read_68d[1] = data_0n[2];
  assign read_68d[2] = data_0n[3];
  assign read_68d[3] = data_0n[4];
  assign read_68d[4] = data_0n[5];
  assign read_68d[5] = data_0n[6];
  assign read_68d[6] = data_0n[7];
  assign read_68d[7] = data_0n[8];
  assign read_68d[8] = data_0n[9];
  assign read_68d[9] = data_0n[10];
  assign read_68d[10] = data_0n[11];
  assign read_68d[11] = data_0n[12];
  assign read_68d[12] = data_0n[13];
  assign read_68d[13] = data_0n[14];
  assign read_68d[14] = data_0n[15];
  assign read_68d[15] = data_0n[16];
  assign read_67d[0] = data_0n[0];
  assign read_67d[1] = data_0n[1];
  assign read_67d[2] = data_0n[2];
  assign read_67d[3] = data_0n[3];
  assign read_67d[4] = data_0n[4];
  assign read_67d[5] = data_0n[5];
  assign read_67d[6] = data_0n[6];
  assign read_67d[7] = data_0n[7];
  assign read_67d[8] = data_0n[8];
  assign read_67d[9] = data_0n[9];
  assign read_67d[10] = data_0n[10];
  assign read_67d[11] = data_0n[11];
  assign read_67d[12] = data_0n[12];
  assign read_67d[13] = data_0n[13];
  assign read_67d[14] = data_0n[14];
  assign read_67d[15] = data_0n[15];
  assign read_67d[16] = data_0n[16];
  assign read_66d[0] = data_0n[0];
  assign read_66d[1] = data_0n[1];
  assign read_66d[2] = data_0n[2];
  assign read_66d[3] = data_0n[3];
  assign read_66d[4] = data_0n[4];
  assign read_66d[5] = data_0n[5];
  assign read_66d[6] = data_0n[6];
  assign read_66d[7] = data_0n[7];
  assign read_66d[8] = data_0n[8];
  assign read_66d[9] = data_0n[9];
  assign read_66d[10] = data_0n[10];
  assign read_66d[11] = data_0n[11];
  assign read_66d[12] = data_0n[12];
  assign read_66d[13] = data_0n[13];
  assign read_66d[14] = data_0n[14];
  assign read_66d[15] = data_0n[15];
  assign read_66d[16] = data_0n[16];
  assign read_65d[0] = data_0n[0];
  assign read_65d[1] = data_0n[1];
  assign read_65d[2] = data_0n[2];
  assign read_65d[3] = data_0n[3];
  assign read_65d[4] = data_0n[4];
  assign read_65d[5] = data_0n[5];
  assign read_65d[6] = data_0n[6];
  assign read_65d[7] = data_0n[7];
  assign read_65d[8] = data_0n[8];
  assign read_65d[9] = data_0n[9];
  assign read_65d[10] = data_0n[10];
  assign read_65d[11] = data_0n[11];
  assign read_65d[12] = data_0n[12];
  assign read_65d[13] = data_0n[13];
  assign read_65d[14] = data_0n[14];
  assign read_65d[15] = data_0n[15];
  assign read_65d[16] = data_0n[16];
  assign read_64d[0] = data_0n[0];
  assign read_64d[1] = data_0n[1];
  assign read_64d[2] = data_0n[2];
  assign read_64d[3] = data_0n[3];
  assign read_64d[4] = data_0n[4];
  assign read_64d[5] = data_0n[5];
  assign read_64d[6] = data_0n[6];
  assign read_64d[7] = data_0n[7];
  assign read_64d[8] = data_0n[8];
  assign read_64d[9] = data_0n[9];
  assign read_64d[10] = data_0n[10];
  assign read_64d[11] = data_0n[11];
  assign read_64d[12] = data_0n[12];
  assign read_64d[13] = data_0n[13];
  assign read_64d[14] = data_0n[14];
  assign read_64d[15] = data_0n[15];
  assign read_64d[16] = data_0n[16];
  assign read_63d = data_0n[0];
  assign read_62d = data_0n[1];
  assign read_61d = data_0n[0];
  assign read_60d = data_0n[1];
  assign read_59d = data_0n[16];
  assign read_58d[0] = data_0n[1];
  assign read_58d[1] = data_0n[2];
  assign read_58d[2] = data_0n[3];
  assign read_58d[3] = data_0n[4];
  assign read_58d[4] = data_0n[5];
  assign read_58d[5] = data_0n[6];
  assign read_58d[6] = data_0n[7];
  assign read_58d[7] = data_0n[8];
  assign read_58d[8] = data_0n[9];
  assign read_58d[9] = data_0n[10];
  assign read_58d[10] = data_0n[11];
  assign read_58d[11] = data_0n[12];
  assign read_58d[12] = data_0n[13];
  assign read_58d[13] = data_0n[14];
  assign read_58d[14] = data_0n[15];
  assign read_58d[15] = data_0n[16];
  assign read_57d[0] = data_0n[0];
  assign read_57d[1] = data_0n[1];
  assign read_57d[2] = data_0n[2];
  assign read_57d[3] = data_0n[3];
  assign read_57d[4] = data_0n[4];
  assign read_57d[5] = data_0n[5];
  assign read_57d[6] = data_0n[6];
  assign read_57d[7] = data_0n[7];
  assign read_57d[8] = data_0n[8];
  assign read_57d[9] = data_0n[9];
  assign read_57d[10] = data_0n[10];
  assign read_57d[11] = data_0n[11];
  assign read_57d[12] = data_0n[12];
  assign read_57d[13] = data_0n[13];
  assign read_57d[14] = data_0n[14];
  assign read_57d[15] = data_0n[15];
  assign read_57d[16] = data_0n[16];
  assign read_56d[0] = data_0n[0];
  assign read_56d[1] = data_0n[1];
  assign read_56d[2] = data_0n[2];
  assign read_56d[3] = data_0n[3];
  assign read_56d[4] = data_0n[4];
  assign read_56d[5] = data_0n[5];
  assign read_56d[6] = data_0n[6];
  assign read_56d[7] = data_0n[7];
  assign read_56d[8] = data_0n[8];
  assign read_56d[9] = data_0n[9];
  assign read_56d[10] = data_0n[10];
  assign read_56d[11] = data_0n[11];
  assign read_56d[12] = data_0n[12];
  assign read_56d[13] = data_0n[13];
  assign read_56d[14] = data_0n[14];
  assign read_56d[15] = data_0n[15];
  assign read_56d[16] = data_0n[16];
  assign read_55d[0] = data_0n[0];
  assign read_55d[1] = data_0n[1];
  assign read_55d[2] = data_0n[2];
  assign read_55d[3] = data_0n[3];
  assign read_55d[4] = data_0n[4];
  assign read_55d[5] = data_0n[5];
  assign read_55d[6] = data_0n[6];
  assign read_55d[7] = data_0n[7];
  assign read_55d[8] = data_0n[8];
  assign read_55d[9] = data_0n[9];
  assign read_55d[10] = data_0n[10];
  assign read_55d[11] = data_0n[11];
  assign read_55d[12] = data_0n[12];
  assign read_55d[13] = data_0n[13];
  assign read_55d[14] = data_0n[14];
  assign read_55d[15] = data_0n[15];
  assign read_55d[16] = data_0n[16];
  assign read_54d[0] = data_0n[0];
  assign read_54d[1] = data_0n[1];
  assign read_54d[2] = data_0n[2];
  assign read_54d[3] = data_0n[3];
  assign read_54d[4] = data_0n[4];
  assign read_54d[5] = data_0n[5];
  assign read_54d[6] = data_0n[6];
  assign read_54d[7] = data_0n[7];
  assign read_54d[8] = data_0n[8];
  assign read_54d[9] = data_0n[9];
  assign read_54d[10] = data_0n[10];
  assign read_54d[11] = data_0n[11];
  assign read_54d[12] = data_0n[12];
  assign read_54d[13] = data_0n[13];
  assign read_54d[14] = data_0n[14];
  assign read_54d[15] = data_0n[15];
  assign read_54d[16] = data_0n[16];
  assign read_53d = data_0n[0];
  assign read_52d = data_0n[1];
  assign read_51d = data_0n[0];
  assign read_50d = data_0n[1];
  assign read_49d = data_0n[16];
  assign read_48d[0] = data_0n[1];
  assign read_48d[1] = data_0n[2];
  assign read_48d[2] = data_0n[3];
  assign read_48d[3] = data_0n[4];
  assign read_48d[4] = data_0n[5];
  assign read_48d[5] = data_0n[6];
  assign read_48d[6] = data_0n[7];
  assign read_48d[7] = data_0n[8];
  assign read_48d[8] = data_0n[9];
  assign read_48d[9] = data_0n[10];
  assign read_48d[10] = data_0n[11];
  assign read_48d[11] = data_0n[12];
  assign read_48d[12] = data_0n[13];
  assign read_48d[13] = data_0n[14];
  assign read_48d[14] = data_0n[15];
  assign read_48d[15] = data_0n[16];
  assign read_47d[0] = data_0n[0];
  assign read_47d[1] = data_0n[1];
  assign read_47d[2] = data_0n[2];
  assign read_47d[3] = data_0n[3];
  assign read_47d[4] = data_0n[4];
  assign read_47d[5] = data_0n[5];
  assign read_47d[6] = data_0n[6];
  assign read_47d[7] = data_0n[7];
  assign read_47d[8] = data_0n[8];
  assign read_47d[9] = data_0n[9];
  assign read_47d[10] = data_0n[10];
  assign read_47d[11] = data_0n[11];
  assign read_47d[12] = data_0n[12];
  assign read_47d[13] = data_0n[13];
  assign read_47d[14] = data_0n[14];
  assign read_47d[15] = data_0n[15];
  assign read_47d[16] = data_0n[16];
  assign read_46d[0] = data_0n[0];
  assign read_46d[1] = data_0n[1];
  assign read_46d[2] = data_0n[2];
  assign read_46d[3] = data_0n[3];
  assign read_46d[4] = data_0n[4];
  assign read_46d[5] = data_0n[5];
  assign read_46d[6] = data_0n[6];
  assign read_46d[7] = data_0n[7];
  assign read_46d[8] = data_0n[8];
  assign read_46d[9] = data_0n[9];
  assign read_46d[10] = data_0n[10];
  assign read_46d[11] = data_0n[11];
  assign read_46d[12] = data_0n[12];
  assign read_46d[13] = data_0n[13];
  assign read_46d[14] = data_0n[14];
  assign read_46d[15] = data_0n[15];
  assign read_46d[16] = data_0n[16];
  assign read_45d[0] = data_0n[0];
  assign read_45d[1] = data_0n[1];
  assign read_45d[2] = data_0n[2];
  assign read_45d[3] = data_0n[3];
  assign read_45d[4] = data_0n[4];
  assign read_45d[5] = data_0n[5];
  assign read_45d[6] = data_0n[6];
  assign read_45d[7] = data_0n[7];
  assign read_45d[8] = data_0n[8];
  assign read_45d[9] = data_0n[9];
  assign read_45d[10] = data_0n[10];
  assign read_45d[11] = data_0n[11];
  assign read_45d[12] = data_0n[12];
  assign read_45d[13] = data_0n[13];
  assign read_45d[14] = data_0n[14];
  assign read_45d[15] = data_0n[15];
  assign read_45d[16] = data_0n[16];
  assign read_44d[0] = data_0n[0];
  assign read_44d[1] = data_0n[1];
  assign read_44d[2] = data_0n[2];
  assign read_44d[3] = data_0n[3];
  assign read_44d[4] = data_0n[4];
  assign read_44d[5] = data_0n[5];
  assign read_44d[6] = data_0n[6];
  assign read_44d[7] = data_0n[7];
  assign read_44d[8] = data_0n[8];
  assign read_44d[9] = data_0n[9];
  assign read_44d[10] = data_0n[10];
  assign read_44d[11] = data_0n[11];
  assign read_44d[12] = data_0n[12];
  assign read_44d[13] = data_0n[13];
  assign read_44d[14] = data_0n[14];
  assign read_44d[15] = data_0n[15];
  assign read_44d[16] = data_0n[16];
  assign read_43d = data_0n[0];
  assign read_42d = data_0n[1];
  assign read_41d = data_0n[0];
  assign read_40d = data_0n[1];
  assign read_39d = data_0n[16];
  assign read_38d[0] = data_0n[1];
  assign read_38d[1] = data_0n[2];
  assign read_38d[2] = data_0n[3];
  assign read_38d[3] = data_0n[4];
  assign read_38d[4] = data_0n[5];
  assign read_38d[5] = data_0n[6];
  assign read_38d[6] = data_0n[7];
  assign read_38d[7] = data_0n[8];
  assign read_38d[8] = data_0n[9];
  assign read_38d[9] = data_0n[10];
  assign read_38d[10] = data_0n[11];
  assign read_38d[11] = data_0n[12];
  assign read_38d[12] = data_0n[13];
  assign read_38d[13] = data_0n[14];
  assign read_38d[14] = data_0n[15];
  assign read_38d[15] = data_0n[16];
  assign read_37d[0] = data_0n[0];
  assign read_37d[1] = data_0n[1];
  assign read_37d[2] = data_0n[2];
  assign read_37d[3] = data_0n[3];
  assign read_37d[4] = data_0n[4];
  assign read_37d[5] = data_0n[5];
  assign read_37d[6] = data_0n[6];
  assign read_37d[7] = data_0n[7];
  assign read_37d[8] = data_0n[8];
  assign read_37d[9] = data_0n[9];
  assign read_37d[10] = data_0n[10];
  assign read_37d[11] = data_0n[11];
  assign read_37d[12] = data_0n[12];
  assign read_37d[13] = data_0n[13];
  assign read_37d[14] = data_0n[14];
  assign read_37d[15] = data_0n[15];
  assign read_37d[16] = data_0n[16];
  assign read_36d[0] = data_0n[0];
  assign read_36d[1] = data_0n[1];
  assign read_36d[2] = data_0n[2];
  assign read_36d[3] = data_0n[3];
  assign read_36d[4] = data_0n[4];
  assign read_36d[5] = data_0n[5];
  assign read_36d[6] = data_0n[6];
  assign read_36d[7] = data_0n[7];
  assign read_36d[8] = data_0n[8];
  assign read_36d[9] = data_0n[9];
  assign read_36d[10] = data_0n[10];
  assign read_36d[11] = data_0n[11];
  assign read_36d[12] = data_0n[12];
  assign read_36d[13] = data_0n[13];
  assign read_36d[14] = data_0n[14];
  assign read_36d[15] = data_0n[15];
  assign read_36d[16] = data_0n[16];
  assign read_35d[0] = data_0n[0];
  assign read_35d[1] = data_0n[1];
  assign read_35d[2] = data_0n[2];
  assign read_35d[3] = data_0n[3];
  assign read_35d[4] = data_0n[4];
  assign read_35d[5] = data_0n[5];
  assign read_35d[6] = data_0n[6];
  assign read_35d[7] = data_0n[7];
  assign read_35d[8] = data_0n[8];
  assign read_35d[9] = data_0n[9];
  assign read_35d[10] = data_0n[10];
  assign read_35d[11] = data_0n[11];
  assign read_35d[12] = data_0n[12];
  assign read_35d[13] = data_0n[13];
  assign read_35d[14] = data_0n[14];
  assign read_35d[15] = data_0n[15];
  assign read_35d[16] = data_0n[16];
  assign read_34d[0] = data_0n[0];
  assign read_34d[1] = data_0n[1];
  assign read_34d[2] = data_0n[2];
  assign read_34d[3] = data_0n[3];
  assign read_34d[4] = data_0n[4];
  assign read_34d[5] = data_0n[5];
  assign read_34d[6] = data_0n[6];
  assign read_34d[7] = data_0n[7];
  assign read_34d[8] = data_0n[8];
  assign read_34d[9] = data_0n[9];
  assign read_34d[10] = data_0n[10];
  assign read_34d[11] = data_0n[11];
  assign read_34d[12] = data_0n[12];
  assign read_34d[13] = data_0n[13];
  assign read_34d[14] = data_0n[14];
  assign read_34d[15] = data_0n[15];
  assign read_34d[16] = data_0n[16];
  assign read_33d = data_0n[0];
  assign read_32d = data_0n[1];
  assign read_31d = data_0n[0];
  assign read_30d = data_0n[1];
  assign read_29d = data_0n[16];
  assign read_28d[0] = data_0n[1];
  assign read_28d[1] = data_0n[2];
  assign read_28d[2] = data_0n[3];
  assign read_28d[3] = data_0n[4];
  assign read_28d[4] = data_0n[5];
  assign read_28d[5] = data_0n[6];
  assign read_28d[6] = data_0n[7];
  assign read_28d[7] = data_0n[8];
  assign read_28d[8] = data_0n[9];
  assign read_28d[9] = data_0n[10];
  assign read_28d[10] = data_0n[11];
  assign read_28d[11] = data_0n[12];
  assign read_28d[12] = data_0n[13];
  assign read_28d[13] = data_0n[14];
  assign read_28d[14] = data_0n[15];
  assign read_28d[15] = data_0n[16];
  assign read_27d[0] = data_0n[0];
  assign read_27d[1] = data_0n[1];
  assign read_27d[2] = data_0n[2];
  assign read_27d[3] = data_0n[3];
  assign read_27d[4] = data_0n[4];
  assign read_27d[5] = data_0n[5];
  assign read_27d[6] = data_0n[6];
  assign read_27d[7] = data_0n[7];
  assign read_27d[8] = data_0n[8];
  assign read_27d[9] = data_0n[9];
  assign read_27d[10] = data_0n[10];
  assign read_27d[11] = data_0n[11];
  assign read_27d[12] = data_0n[12];
  assign read_27d[13] = data_0n[13];
  assign read_27d[14] = data_0n[14];
  assign read_27d[15] = data_0n[15];
  assign read_27d[16] = data_0n[16];
  assign read_26d[0] = data_0n[0];
  assign read_26d[1] = data_0n[1];
  assign read_26d[2] = data_0n[2];
  assign read_26d[3] = data_0n[3];
  assign read_26d[4] = data_0n[4];
  assign read_26d[5] = data_0n[5];
  assign read_26d[6] = data_0n[6];
  assign read_26d[7] = data_0n[7];
  assign read_26d[8] = data_0n[8];
  assign read_26d[9] = data_0n[9];
  assign read_26d[10] = data_0n[10];
  assign read_26d[11] = data_0n[11];
  assign read_26d[12] = data_0n[12];
  assign read_26d[13] = data_0n[13];
  assign read_26d[14] = data_0n[14];
  assign read_26d[15] = data_0n[15];
  assign read_26d[16] = data_0n[16];
  assign read_25d[0] = data_0n[0];
  assign read_25d[1] = data_0n[1];
  assign read_25d[2] = data_0n[2];
  assign read_25d[3] = data_0n[3];
  assign read_25d[4] = data_0n[4];
  assign read_25d[5] = data_0n[5];
  assign read_25d[6] = data_0n[6];
  assign read_25d[7] = data_0n[7];
  assign read_25d[8] = data_0n[8];
  assign read_25d[9] = data_0n[9];
  assign read_25d[10] = data_0n[10];
  assign read_25d[11] = data_0n[11];
  assign read_25d[12] = data_0n[12];
  assign read_25d[13] = data_0n[13];
  assign read_25d[14] = data_0n[14];
  assign read_25d[15] = data_0n[15];
  assign read_25d[16] = data_0n[16];
  assign read_24d[0] = data_0n[0];
  assign read_24d[1] = data_0n[1];
  assign read_24d[2] = data_0n[2];
  assign read_24d[3] = data_0n[3];
  assign read_24d[4] = data_0n[4];
  assign read_24d[5] = data_0n[5];
  assign read_24d[6] = data_0n[6];
  assign read_24d[7] = data_0n[7];
  assign read_24d[8] = data_0n[8];
  assign read_24d[9] = data_0n[9];
  assign read_24d[10] = data_0n[10];
  assign read_24d[11] = data_0n[11];
  assign read_24d[12] = data_0n[12];
  assign read_24d[13] = data_0n[13];
  assign read_24d[14] = data_0n[14];
  assign read_24d[15] = data_0n[15];
  assign read_24d[16] = data_0n[16];
  assign read_23d = data_0n[0];
  assign read_22d = data_0n[1];
  assign read_21d = data_0n[0];
  assign read_20d = data_0n[1];
  assign read_19d = data_0n[16];
  assign read_18d[0] = data_0n[1];
  assign read_18d[1] = data_0n[2];
  assign read_18d[2] = data_0n[3];
  assign read_18d[3] = data_0n[4];
  assign read_18d[4] = data_0n[5];
  assign read_18d[5] = data_0n[6];
  assign read_18d[6] = data_0n[7];
  assign read_18d[7] = data_0n[8];
  assign read_18d[8] = data_0n[9];
  assign read_18d[9] = data_0n[10];
  assign read_18d[10] = data_0n[11];
  assign read_18d[11] = data_0n[12];
  assign read_18d[12] = data_0n[13];
  assign read_18d[13] = data_0n[14];
  assign read_18d[14] = data_0n[15];
  assign read_18d[15] = data_0n[16];
  assign read_17d[0] = data_0n[0];
  assign read_17d[1] = data_0n[1];
  assign read_17d[2] = data_0n[2];
  assign read_17d[3] = data_0n[3];
  assign read_17d[4] = data_0n[4];
  assign read_17d[5] = data_0n[5];
  assign read_17d[6] = data_0n[6];
  assign read_17d[7] = data_0n[7];
  assign read_17d[8] = data_0n[8];
  assign read_17d[9] = data_0n[9];
  assign read_17d[10] = data_0n[10];
  assign read_17d[11] = data_0n[11];
  assign read_17d[12] = data_0n[12];
  assign read_17d[13] = data_0n[13];
  assign read_17d[14] = data_0n[14];
  assign read_17d[15] = data_0n[15];
  assign read_17d[16] = data_0n[16];
  assign read_16d[0] = data_0n[0];
  assign read_16d[1] = data_0n[1];
  assign read_16d[2] = data_0n[2];
  assign read_16d[3] = data_0n[3];
  assign read_16d[4] = data_0n[4];
  assign read_16d[5] = data_0n[5];
  assign read_16d[6] = data_0n[6];
  assign read_16d[7] = data_0n[7];
  assign read_16d[8] = data_0n[8];
  assign read_16d[9] = data_0n[9];
  assign read_16d[10] = data_0n[10];
  assign read_16d[11] = data_0n[11];
  assign read_16d[12] = data_0n[12];
  assign read_16d[13] = data_0n[13];
  assign read_16d[14] = data_0n[14];
  assign read_16d[15] = data_0n[15];
  assign read_16d[16] = data_0n[16];
  assign read_15d[0] = data_0n[0];
  assign read_15d[1] = data_0n[1];
  assign read_15d[2] = data_0n[2];
  assign read_15d[3] = data_0n[3];
  assign read_15d[4] = data_0n[4];
  assign read_15d[5] = data_0n[5];
  assign read_15d[6] = data_0n[6];
  assign read_15d[7] = data_0n[7];
  assign read_15d[8] = data_0n[8];
  assign read_15d[9] = data_0n[9];
  assign read_15d[10] = data_0n[10];
  assign read_15d[11] = data_0n[11];
  assign read_15d[12] = data_0n[12];
  assign read_15d[13] = data_0n[13];
  assign read_15d[14] = data_0n[14];
  assign read_15d[15] = data_0n[15];
  assign read_15d[16] = data_0n[16];
  assign read_14d[0] = data_0n[0];
  assign read_14d[1] = data_0n[1];
  assign read_14d[2] = data_0n[2];
  assign read_14d[3] = data_0n[3];
  assign read_14d[4] = data_0n[4];
  assign read_14d[5] = data_0n[5];
  assign read_14d[6] = data_0n[6];
  assign read_14d[7] = data_0n[7];
  assign read_14d[8] = data_0n[8];
  assign read_14d[9] = data_0n[9];
  assign read_14d[10] = data_0n[10];
  assign read_14d[11] = data_0n[11];
  assign read_14d[12] = data_0n[12];
  assign read_14d[13] = data_0n[13];
  assign read_14d[14] = data_0n[14];
  assign read_14d[15] = data_0n[15];
  assign read_14d[16] = data_0n[16];
  assign read_13d = data_0n[0];
  assign read_12d = data_0n[1];
  assign read_11d = data_0n[0];
  assign read_10d = data_0n[1];
  assign read_9d = data_0n[16];
  assign read_8d[0] = data_0n[1];
  assign read_8d[1] = data_0n[2];
  assign read_8d[2] = data_0n[3];
  assign read_8d[3] = data_0n[4];
  assign read_8d[4] = data_0n[5];
  assign read_8d[5] = data_0n[6];
  assign read_8d[6] = data_0n[7];
  assign read_8d[7] = data_0n[8];
  assign read_8d[8] = data_0n[9];
  assign read_8d[9] = data_0n[10];
  assign read_8d[10] = data_0n[11];
  assign read_8d[11] = data_0n[12];
  assign read_8d[12] = data_0n[13];
  assign read_8d[13] = data_0n[14];
  assign read_8d[14] = data_0n[15];
  assign read_8d[15] = data_0n[16];
  assign read_7d[0] = data_0n[0];
  assign read_7d[1] = data_0n[1];
  assign read_7d[2] = data_0n[2];
  assign read_7d[3] = data_0n[3];
  assign read_7d[4] = data_0n[4];
  assign read_7d[5] = data_0n[5];
  assign read_7d[6] = data_0n[6];
  assign read_7d[7] = data_0n[7];
  assign read_7d[8] = data_0n[8];
  assign read_7d[9] = data_0n[9];
  assign read_7d[10] = data_0n[10];
  assign read_7d[11] = data_0n[11];
  assign read_7d[12] = data_0n[12];
  assign read_7d[13] = data_0n[13];
  assign read_7d[14] = data_0n[14];
  assign read_7d[15] = data_0n[15];
  assign read_7d[16] = data_0n[16];
  assign read_6d[0] = data_0n[0];
  assign read_6d[1] = data_0n[1];
  assign read_6d[2] = data_0n[2];
  assign read_6d[3] = data_0n[3];
  assign read_6d[4] = data_0n[4];
  assign read_6d[5] = data_0n[5];
  assign read_6d[6] = data_0n[6];
  assign read_6d[7] = data_0n[7];
  assign read_6d[8] = data_0n[8];
  assign read_6d[9] = data_0n[9];
  assign read_6d[10] = data_0n[10];
  assign read_6d[11] = data_0n[11];
  assign read_6d[12] = data_0n[12];
  assign read_6d[13] = data_0n[13];
  assign read_6d[14] = data_0n[14];
  assign read_6d[15] = data_0n[15];
  assign read_6d[16] = data_0n[16];
  assign read_5d[0] = data_0n[0];
  assign read_5d[1] = data_0n[1];
  assign read_5d[2] = data_0n[2];
  assign read_5d[3] = data_0n[3];
  assign read_5d[4] = data_0n[4];
  assign read_5d[5] = data_0n[5];
  assign read_5d[6] = data_0n[6];
  assign read_5d[7] = data_0n[7];
  assign read_5d[8] = data_0n[8];
  assign read_5d[9] = data_0n[9];
  assign read_5d[10] = data_0n[10];
  assign read_5d[11] = data_0n[11];
  assign read_5d[12] = data_0n[12];
  assign read_5d[13] = data_0n[13];
  assign read_5d[14] = data_0n[14];
  assign read_5d[15] = data_0n[15];
  assign read_5d[16] = data_0n[16];
  assign read_4d[0] = data_0n[0];
  assign read_4d[1] = data_0n[1];
  assign read_4d[2] = data_0n[2];
  assign read_4d[3] = data_0n[3];
  assign read_4d[4] = data_0n[4];
  assign read_4d[5] = data_0n[5];
  assign read_4d[6] = data_0n[6];
  assign read_4d[7] = data_0n[7];
  assign read_4d[8] = data_0n[8];
  assign read_4d[9] = data_0n[9];
  assign read_4d[10] = data_0n[10];
  assign read_4d[11] = data_0n[11];
  assign read_4d[12] = data_0n[12];
  assign read_4d[13] = data_0n[13];
  assign read_4d[14] = data_0n[14];
  assign read_4d[15] = data_0n[15];
  assign read_4d[16] = data_0n[16];
  assign read_3d = data_0n[0];
  assign read_2d = data_0n[1];
  assign read_1d = data_0n[0];
  assign read_0d = data_0n[1];
  LD1 I809 (write_0d[0], bWriteReq_0n, data_0n[0]);
  LD1 I810 (write_0d[1], bWriteReq_0n, data_0n[1]);
  LD1 I811 (write_0d[2], bWriteReq_0n, data_0n[2]);
  LD1 I812 (write_0d[3], bWriteReq_0n, data_0n[3]);
  LD1 I813 (write_0d[4], bWriteReq_0n, data_0n[4]);
  LD1 I814 (write_0d[5], bWriteReq_0n, data_0n[5]);
  LD1 I815 (write_0d[6], bWriteReq_0n, data_0n[6]);
  LD1 I816 (write_0d[7], bWriteReq_0n, data_0n[7]);
  LD1 I817 (write_0d[8], bWriteReq_0n, data_0n[8]);
  LD1 I818 (write_0d[9], bWriteReq_0n, data_0n[9]);
  LD1 I819 (write_0d[10], bWriteReq_0n, data_0n[10]);
  LD1 I820 (write_0d[11], bWriteReq_0n, data_0n[11]);
  LD1 I821 (write_0d[12], bWriteReq_0n, data_0n[12]);
  LD1 I822 (write_0d[13], bWriteReq_0n, data_0n[13]);
  LD1 I823 (write_0d[14], bWriteReq_0n, data_0n[14]);
  LD1 I824 (write_0d[15], bWriteReq_0n, data_0n[15]);
  LD1 I825 (write_0d[16], bWriteReq_0n, data_0n[16]);
  IV I826 (write_0a, nbWriteReq_0n);
  IV I827 (nbWriteReq_0n, bWriteReq_0n);
  IV I828 (bWriteReq_0n, nWriteReq_0n);
  IV I829 (nWriteReq_0n, write_0r);
endmodule

module Balsa_booth__mul8 (
  activate_0r, activate_0a,
  x_0r, x_0a, x_0d,
  y_0r, y_0a, y_0d,
  z_0r, z_0a, z_0d
);
  input activate_0r;
  output activate_0a;
  output x_0r;
  input x_0a;
  input [7:0] x_0d;
  output y_0r;
  input y_0a;
  input [7:0] y_0d;
  output z_0r;
  input z_0a;
  output [15:0] z_0d;
  wire c463_r;
  wire c463_a;
  wire [16:0] c463_d;
  wire c462_r;
  wire c462_a;
  wire c461_r;
  wire c461_a;
  wire c460_r;
  wire c460_a;
  wire c459_r;
  wire c459_a;
  wire [7:0] c459_d;
  wire c458_r;
  wire c458_a;
  wire c457_r;
  wire c457_a;
  wire [7:0] c457_d;
  wire c456_r;
  wire c456_a;
  wire c455_r;
  wire c455_a;
  wire c454_r;
  wire c454_a;
  wire [16:0] c454_d;
  wire c453_r;
  wire c453_a;
  wire [16:0] c453_d;
  wire c452_r;
  wire c452_a;
  wire [8:0] c452_d;
  wire c451_r;
  wire c451_a;
  wire [7:0] c451_d;
  wire c450_r;
  wire c450_a;
  wire c449_r;
  wire c449_a;
  wire [16:0] c449_d;
  wire c448_r;
  wire c448_a;
  wire [16:0] c448_d;
  wire c447_r;
  wire c447_a;
  wire [8:0] c447_d;
  wire c446_r;
  wire c446_a;
  wire [7:0] c446_d;
  wire c445_r;
  wire c445_a;
  wire [7:0] c445_d;
  wire c444_r;
  wire c444_a;
  wire c443_r;
  wire c443_a;
  wire [16:0] c443_d;
  wire c442_r;
  wire c442_a;
  wire [16:0] c442_d;
  wire c441_r;
  wire c441_a;
  wire [8:0] c441_d;
  wire c440_r;
  wire c440_a;
  wire c440_d;
  wire c439_r;
  wire c439_a;
  wire [7:0] c439_d;
  wire c438_r;
  wire c438_a;
  wire c438_d;
  wire c437_r;
  wire c437_a;
  wire c437_d;
  wire c436_r;
  wire c436_a;
  wire c435_r;
  wire c435_a;
  wire c434_r;
  wire c434_a;
  wire c434_d;
  wire c433_r;
  wire c433_a;
  wire c432_r;
  wire c432_a;
  wire c432_d;
  wire c431_r;
  wire c431_a;
  wire c431_d;
  wire c430_r;
  wire c430_a;
  wire c430_d;
  wire c429_r;
  wire c429_a;
  wire c429_d;
  wire c428_r;
  wire c428_a;
  wire c428_d;
  wire c427_r;
  wire c427_a;
  wire [16:0] c427_d;
  wire c426_r;
  wire c426_a;
  wire [16:0] c426_d;
  wire c425_r;
  wire c425_a;
  wire c424_r;
  wire c424_a;
  wire c423_r;
  wire c423_a;
  wire c422_r;
  wire c422_a;
  wire [16:0] c422_d;
  wire c421_r;
  wire c421_a;
  wire [16:0] c421_d;
  wire c420_r;
  wire c420_a;
  wire [15:0] c420_d;
  wire c419_r;
  wire c419_a;
  wire [17:0] c419_d;
  wire c418_r;
  wire c418_a;
  wire [16:0] c418_d;
  wire c417_r;
  wire c417_a;
  wire [16:0] c417_d;
  wire c416_r;
  wire c416_a;
  wire c416_d;
  wire c415_r;
  wire c415_a;
  wire [17:0] c415_d;
  wire c414_r;
  wire c414_a;
  wire [16:0] c414_d;
  wire c413_r;
  wire c413_a;
  wire [16:0] c413_d;
  wire c412_r;
  wire c412_a;
  wire c412_d;
  wire c411_r;
  wire c411_a;
  wire c411_d;
  wire c410_r;
  wire c410_a;
  wire c410_d;
  wire c409_r;
  wire c409_a;
  wire c409_d;
  wire c408_r;
  wire c408_a;
  wire [16:0] c408_d;
  wire c407_r;
  wire c407_a;
  wire [16:0] c407_d;
  wire c406_r;
  wire c406_a;
  wire c405_r;
  wire c405_a;
  wire c404_r;
  wire c404_a;
  wire c403_r;
  wire c403_a;
  wire [16:0] c403_d;
  wire c402_r;
  wire c402_a;
  wire [16:0] c402_d;
  wire c401_r;
  wire c401_a;
  wire [15:0] c401_d;
  wire c400_r;
  wire c400_a;
  wire [17:0] c400_d;
  wire c399_r;
  wire c399_a;
  wire [16:0] c399_d;
  wire c398_r;
  wire c398_a;
  wire [16:0] c398_d;
  wire c397_r;
  wire c397_a;
  wire c397_d;
  wire c396_r;
  wire c396_a;
  wire [17:0] c396_d;
  wire c395_r;
  wire c395_a;
  wire [16:0] c395_d;
  wire c394_r;
  wire c394_a;
  wire [16:0] c394_d;
  wire c393_r;
  wire c393_a;
  wire [16:0] c393_d;
  wire c392_r;
  wire c392_a;
  wire [16:0] c392_d;
  wire c391_r;
  wire c391_a;
  wire c390_r;
  wire c390_a;
  wire c389_r;
  wire c389_a;
  wire c388_r;
  wire c388_a;
  wire [16:0] c388_d;
  wire c387_r;
  wire c387_a;
  wire [16:0] c387_d;
  wire c386_r;
  wire c386_a;
  wire [15:0] c386_d;
  wire c385_r;
  wire c385_a;
  wire c385_d;
  wire c384_r;
  wire c384_a;
  wire c384_d;
  wire c383_r;
  wire c383_a;
  wire c383_d;
  wire c382_r;
  wire c382_a;
  wire c381_r;
  wire c381_a;
  wire c380_r;
  wire c380_a;
  wire c380_d;
  wire c379_r;
  wire c379_a;
  wire c378_r;
  wire c378_a;
  wire c378_d;
  wire c377_r;
  wire c377_a;
  wire c377_d;
  wire c376_r;
  wire c376_a;
  wire c376_d;
  wire c375_r;
  wire c375_a;
  wire c375_d;
  wire c374_r;
  wire c374_a;
  wire c374_d;
  wire c373_r;
  wire c373_a;
  wire [16:0] c373_d;
  wire c372_r;
  wire c372_a;
  wire [16:0] c372_d;
  wire c371_r;
  wire c371_a;
  wire c370_r;
  wire c370_a;
  wire c369_r;
  wire c369_a;
  wire c368_r;
  wire c368_a;
  wire [16:0] c368_d;
  wire c367_r;
  wire c367_a;
  wire [16:0] c367_d;
  wire c366_r;
  wire c366_a;
  wire [15:0] c366_d;
  wire c365_r;
  wire c365_a;
  wire [17:0] c365_d;
  wire c364_r;
  wire c364_a;
  wire [16:0] c364_d;
  wire c363_r;
  wire c363_a;
  wire [16:0] c363_d;
  wire c362_r;
  wire c362_a;
  wire c362_d;
  wire c361_r;
  wire c361_a;
  wire [17:0] c361_d;
  wire c360_r;
  wire c360_a;
  wire [16:0] c360_d;
  wire c359_r;
  wire c359_a;
  wire [16:0] c359_d;
  wire c358_r;
  wire c358_a;
  wire c358_d;
  wire c357_r;
  wire c357_a;
  wire c357_d;
  wire c356_r;
  wire c356_a;
  wire c356_d;
  wire c355_r;
  wire c355_a;
  wire c355_d;
  wire c354_r;
  wire c354_a;
  wire [16:0] c354_d;
  wire c353_r;
  wire c353_a;
  wire [16:0] c353_d;
  wire c352_r;
  wire c352_a;
  wire c351_r;
  wire c351_a;
  wire c350_r;
  wire c350_a;
  wire c349_r;
  wire c349_a;
  wire [16:0] c349_d;
  wire c348_r;
  wire c348_a;
  wire [16:0] c348_d;
  wire c347_r;
  wire c347_a;
  wire [15:0] c347_d;
  wire c346_r;
  wire c346_a;
  wire [17:0] c346_d;
  wire c345_r;
  wire c345_a;
  wire [16:0] c345_d;
  wire c344_r;
  wire c344_a;
  wire [16:0] c344_d;
  wire c343_r;
  wire c343_a;
  wire c343_d;
  wire c342_r;
  wire c342_a;
  wire [17:0] c342_d;
  wire c341_r;
  wire c341_a;
  wire [16:0] c341_d;
  wire c340_r;
  wire c340_a;
  wire [16:0] c340_d;
  wire c339_r;
  wire c339_a;
  wire [16:0] c339_d;
  wire c338_r;
  wire c338_a;
  wire [16:0] c338_d;
  wire c337_r;
  wire c337_a;
  wire c336_r;
  wire c336_a;
  wire c335_r;
  wire c335_a;
  wire c334_r;
  wire c334_a;
  wire [16:0] c334_d;
  wire c333_r;
  wire c333_a;
  wire [16:0] c333_d;
  wire c332_r;
  wire c332_a;
  wire [15:0] c332_d;
  wire c331_r;
  wire c331_a;
  wire c331_d;
  wire c330_r;
  wire c330_a;
  wire c330_d;
  wire c329_r;
  wire c329_a;
  wire c329_d;
  wire c328_r;
  wire c328_a;
  wire c327_r;
  wire c327_a;
  wire c326_r;
  wire c326_a;
  wire c326_d;
  wire c325_r;
  wire c325_a;
  wire c324_r;
  wire c324_a;
  wire c324_d;
  wire c323_r;
  wire c323_a;
  wire c323_d;
  wire c322_r;
  wire c322_a;
  wire c322_d;
  wire c321_r;
  wire c321_a;
  wire c321_d;
  wire c320_r;
  wire c320_a;
  wire c320_d;
  wire c319_r;
  wire c319_a;
  wire [16:0] c319_d;
  wire c318_r;
  wire c318_a;
  wire [16:0] c318_d;
  wire c317_r;
  wire c317_a;
  wire c316_r;
  wire c316_a;
  wire c315_r;
  wire c315_a;
  wire c314_r;
  wire c314_a;
  wire [16:0] c314_d;
  wire c313_r;
  wire c313_a;
  wire [16:0] c313_d;
  wire c312_r;
  wire c312_a;
  wire [15:0] c312_d;
  wire c311_r;
  wire c311_a;
  wire [17:0] c311_d;
  wire c310_r;
  wire c310_a;
  wire [16:0] c310_d;
  wire c309_r;
  wire c309_a;
  wire [16:0] c309_d;
  wire c308_r;
  wire c308_a;
  wire c308_d;
  wire c307_r;
  wire c307_a;
  wire [17:0] c307_d;
  wire c306_r;
  wire c306_a;
  wire [16:0] c306_d;
  wire c305_r;
  wire c305_a;
  wire [16:0] c305_d;
  wire c304_r;
  wire c304_a;
  wire c304_d;
  wire c303_r;
  wire c303_a;
  wire c303_d;
  wire c302_r;
  wire c302_a;
  wire c302_d;
  wire c301_r;
  wire c301_a;
  wire c301_d;
  wire c300_r;
  wire c300_a;
  wire [16:0] c300_d;
  wire c299_r;
  wire c299_a;
  wire [16:0] c299_d;
  wire c298_r;
  wire c298_a;
  wire c297_r;
  wire c297_a;
  wire c296_r;
  wire c296_a;
  wire c295_r;
  wire c295_a;
  wire [16:0] c295_d;
  wire c294_r;
  wire c294_a;
  wire [16:0] c294_d;
  wire c293_r;
  wire c293_a;
  wire [15:0] c293_d;
  wire c292_r;
  wire c292_a;
  wire [17:0] c292_d;
  wire c291_r;
  wire c291_a;
  wire [16:0] c291_d;
  wire c290_r;
  wire c290_a;
  wire [16:0] c290_d;
  wire c289_r;
  wire c289_a;
  wire c289_d;
  wire c288_r;
  wire c288_a;
  wire [17:0] c288_d;
  wire c287_r;
  wire c287_a;
  wire [16:0] c287_d;
  wire c286_r;
  wire c286_a;
  wire [16:0] c286_d;
  wire c285_r;
  wire c285_a;
  wire [16:0] c285_d;
  wire c284_r;
  wire c284_a;
  wire [16:0] c284_d;
  wire c283_r;
  wire c283_a;
  wire c282_r;
  wire c282_a;
  wire c281_r;
  wire c281_a;
  wire c280_r;
  wire c280_a;
  wire [16:0] c280_d;
  wire c279_r;
  wire c279_a;
  wire [16:0] c279_d;
  wire c278_r;
  wire c278_a;
  wire [15:0] c278_d;
  wire c277_r;
  wire c277_a;
  wire c277_d;
  wire c276_r;
  wire c276_a;
  wire c276_d;
  wire c275_r;
  wire c275_a;
  wire c275_d;
  wire c274_r;
  wire c274_a;
  wire c273_r;
  wire c273_a;
  wire c272_r;
  wire c272_a;
  wire c272_d;
  wire c271_r;
  wire c271_a;
  wire c270_r;
  wire c270_a;
  wire c270_d;
  wire c269_r;
  wire c269_a;
  wire c269_d;
  wire c268_r;
  wire c268_a;
  wire c268_d;
  wire c267_r;
  wire c267_a;
  wire c267_d;
  wire c266_r;
  wire c266_a;
  wire c266_d;
  wire c265_r;
  wire c265_a;
  wire [16:0] c265_d;
  wire c264_r;
  wire c264_a;
  wire [16:0] c264_d;
  wire c263_r;
  wire c263_a;
  wire c262_r;
  wire c262_a;
  wire c261_r;
  wire c261_a;
  wire c260_r;
  wire c260_a;
  wire [16:0] c260_d;
  wire c259_r;
  wire c259_a;
  wire [16:0] c259_d;
  wire c258_r;
  wire c258_a;
  wire [15:0] c258_d;
  wire c257_r;
  wire c257_a;
  wire [17:0] c257_d;
  wire c256_r;
  wire c256_a;
  wire [16:0] c256_d;
  wire c255_r;
  wire c255_a;
  wire [16:0] c255_d;
  wire c254_r;
  wire c254_a;
  wire c254_d;
  wire c253_r;
  wire c253_a;
  wire [17:0] c253_d;
  wire c252_r;
  wire c252_a;
  wire [16:0] c252_d;
  wire c251_r;
  wire c251_a;
  wire [16:0] c251_d;
  wire c250_r;
  wire c250_a;
  wire c250_d;
  wire c249_r;
  wire c249_a;
  wire c249_d;
  wire c248_r;
  wire c248_a;
  wire c248_d;
  wire c247_r;
  wire c247_a;
  wire c247_d;
  wire c246_r;
  wire c246_a;
  wire [16:0] c246_d;
  wire c245_r;
  wire c245_a;
  wire [16:0] c245_d;
  wire c244_r;
  wire c244_a;
  wire c243_r;
  wire c243_a;
  wire c242_r;
  wire c242_a;
  wire c241_r;
  wire c241_a;
  wire [16:0] c241_d;
  wire c240_r;
  wire c240_a;
  wire [16:0] c240_d;
  wire c239_r;
  wire c239_a;
  wire [15:0] c239_d;
  wire c238_r;
  wire c238_a;
  wire [17:0] c238_d;
  wire c237_r;
  wire c237_a;
  wire [16:0] c237_d;
  wire c236_r;
  wire c236_a;
  wire [16:0] c236_d;
  wire c235_r;
  wire c235_a;
  wire c235_d;
  wire c234_r;
  wire c234_a;
  wire [17:0] c234_d;
  wire c233_r;
  wire c233_a;
  wire [16:0] c233_d;
  wire c232_r;
  wire c232_a;
  wire [16:0] c232_d;
  wire c231_r;
  wire c231_a;
  wire [16:0] c231_d;
  wire c230_r;
  wire c230_a;
  wire [16:0] c230_d;
  wire c229_r;
  wire c229_a;
  wire c228_r;
  wire c228_a;
  wire c227_r;
  wire c227_a;
  wire c226_r;
  wire c226_a;
  wire [16:0] c226_d;
  wire c225_r;
  wire c225_a;
  wire [16:0] c225_d;
  wire c224_r;
  wire c224_a;
  wire [15:0] c224_d;
  wire c223_r;
  wire c223_a;
  wire c223_d;
  wire c222_r;
  wire c222_a;
  wire c222_d;
  wire c221_r;
  wire c221_a;
  wire c221_d;
  wire c220_r;
  wire c220_a;
  wire c219_r;
  wire c219_a;
  wire c218_r;
  wire c218_a;
  wire c218_d;
  wire c217_r;
  wire c217_a;
  wire c216_r;
  wire c216_a;
  wire c216_d;
  wire c215_r;
  wire c215_a;
  wire c215_d;
  wire c214_r;
  wire c214_a;
  wire c214_d;
  wire c213_r;
  wire c213_a;
  wire c213_d;
  wire c212_r;
  wire c212_a;
  wire c212_d;
  wire c211_r;
  wire c211_a;
  wire [16:0] c211_d;
  wire c210_r;
  wire c210_a;
  wire [16:0] c210_d;
  wire c209_r;
  wire c209_a;
  wire c208_r;
  wire c208_a;
  wire c207_r;
  wire c207_a;
  wire c206_r;
  wire c206_a;
  wire [16:0] c206_d;
  wire c205_r;
  wire c205_a;
  wire [16:0] c205_d;
  wire c204_r;
  wire c204_a;
  wire [15:0] c204_d;
  wire c203_r;
  wire c203_a;
  wire [17:0] c203_d;
  wire c202_r;
  wire c202_a;
  wire [16:0] c202_d;
  wire c201_r;
  wire c201_a;
  wire [16:0] c201_d;
  wire c200_r;
  wire c200_a;
  wire c200_d;
  wire c199_r;
  wire c199_a;
  wire [17:0] c199_d;
  wire c198_r;
  wire c198_a;
  wire [16:0] c198_d;
  wire c197_r;
  wire c197_a;
  wire [16:0] c197_d;
  wire c196_r;
  wire c196_a;
  wire c196_d;
  wire c195_r;
  wire c195_a;
  wire c195_d;
  wire c194_r;
  wire c194_a;
  wire c194_d;
  wire c193_r;
  wire c193_a;
  wire c193_d;
  wire c192_r;
  wire c192_a;
  wire [16:0] c192_d;
  wire c191_r;
  wire c191_a;
  wire [16:0] c191_d;
  wire c190_r;
  wire c190_a;
  wire c189_r;
  wire c189_a;
  wire c188_r;
  wire c188_a;
  wire c187_r;
  wire c187_a;
  wire [16:0] c187_d;
  wire c186_r;
  wire c186_a;
  wire [16:0] c186_d;
  wire c185_r;
  wire c185_a;
  wire [15:0] c185_d;
  wire c184_r;
  wire c184_a;
  wire [17:0] c184_d;
  wire c183_r;
  wire c183_a;
  wire [16:0] c183_d;
  wire c182_r;
  wire c182_a;
  wire [16:0] c182_d;
  wire c181_r;
  wire c181_a;
  wire c181_d;
  wire c180_r;
  wire c180_a;
  wire [17:0] c180_d;
  wire c179_r;
  wire c179_a;
  wire [16:0] c179_d;
  wire c178_r;
  wire c178_a;
  wire [16:0] c178_d;
  wire c177_r;
  wire c177_a;
  wire [16:0] c177_d;
  wire c176_r;
  wire c176_a;
  wire [16:0] c176_d;
  wire c175_r;
  wire c175_a;
  wire c174_r;
  wire c174_a;
  wire c173_r;
  wire c173_a;
  wire c172_r;
  wire c172_a;
  wire [16:0] c172_d;
  wire c171_r;
  wire c171_a;
  wire [16:0] c171_d;
  wire c170_r;
  wire c170_a;
  wire [15:0] c170_d;
  wire c169_r;
  wire c169_a;
  wire c169_d;
  wire c168_r;
  wire c168_a;
  wire c168_d;
  wire c167_r;
  wire c167_a;
  wire c167_d;
  wire c166_r;
  wire c166_a;
  wire c165_r;
  wire c165_a;
  wire c164_r;
  wire c164_a;
  wire c164_d;
  wire c163_r;
  wire c163_a;
  wire c162_r;
  wire c162_a;
  wire c162_d;
  wire c161_r;
  wire c161_a;
  wire c161_d;
  wire c160_r;
  wire c160_a;
  wire c160_d;
  wire c159_r;
  wire c159_a;
  wire c159_d;
  wire c158_r;
  wire c158_a;
  wire c158_d;
  wire c157_r;
  wire c157_a;
  wire [16:0] c157_d;
  wire c156_r;
  wire c156_a;
  wire [16:0] c156_d;
  wire c155_r;
  wire c155_a;
  wire c154_r;
  wire c154_a;
  wire c153_r;
  wire c153_a;
  wire c152_r;
  wire c152_a;
  wire [16:0] c152_d;
  wire c151_r;
  wire c151_a;
  wire [16:0] c151_d;
  wire c150_r;
  wire c150_a;
  wire [15:0] c150_d;
  wire c149_r;
  wire c149_a;
  wire [17:0] c149_d;
  wire c148_r;
  wire c148_a;
  wire [16:0] c148_d;
  wire c147_r;
  wire c147_a;
  wire [16:0] c147_d;
  wire c146_r;
  wire c146_a;
  wire c146_d;
  wire c145_r;
  wire c145_a;
  wire [17:0] c145_d;
  wire c144_r;
  wire c144_a;
  wire [16:0] c144_d;
  wire c143_r;
  wire c143_a;
  wire [16:0] c143_d;
  wire c142_r;
  wire c142_a;
  wire c142_d;
  wire c141_r;
  wire c141_a;
  wire c141_d;
  wire c140_r;
  wire c140_a;
  wire c140_d;
  wire c139_r;
  wire c139_a;
  wire c139_d;
  wire c138_r;
  wire c138_a;
  wire [16:0] c138_d;
  wire c137_r;
  wire c137_a;
  wire [16:0] c137_d;
  wire c136_r;
  wire c136_a;
  wire c135_r;
  wire c135_a;
  wire c134_r;
  wire c134_a;
  wire c133_r;
  wire c133_a;
  wire [16:0] c133_d;
  wire c132_r;
  wire c132_a;
  wire [16:0] c132_d;
  wire c131_r;
  wire c131_a;
  wire [15:0] c131_d;
  wire c130_r;
  wire c130_a;
  wire [17:0] c130_d;
  wire c129_r;
  wire c129_a;
  wire [16:0] c129_d;
  wire c128_r;
  wire c128_a;
  wire [16:0] c128_d;
  wire c127_r;
  wire c127_a;
  wire c127_d;
  wire c126_r;
  wire c126_a;
  wire [17:0] c126_d;
  wire c125_r;
  wire c125_a;
  wire [16:0] c125_d;
  wire c124_r;
  wire c124_a;
  wire [16:0] c124_d;
  wire c123_r;
  wire c123_a;
  wire [16:0] c123_d;
  wire c122_r;
  wire c122_a;
  wire [16:0] c122_d;
  wire c121_r;
  wire c121_a;
  wire c120_r;
  wire c120_a;
  wire c119_r;
  wire c119_a;
  wire c118_r;
  wire c118_a;
  wire [16:0] c118_d;
  wire c117_r;
  wire c117_a;
  wire [16:0] c117_d;
  wire c116_r;
  wire c116_a;
  wire [15:0] c116_d;
  wire c115_r;
  wire c115_a;
  wire c115_d;
  wire c114_r;
  wire c114_a;
  wire c114_d;
  wire c113_r;
  wire c113_a;
  wire c113_d;
  wire c112_r;
  wire c112_a;
  wire c111_r;
  wire c111_a;
  wire c110_r;
  wire c110_a;
  wire c110_d;
  wire c109_r;
  wire c109_a;
  wire c108_r;
  wire c108_a;
  wire c108_d;
  wire c107_r;
  wire c107_a;
  wire c107_d;
  wire c106_r;
  wire c106_a;
  wire c106_d;
  wire c105_r;
  wire c105_a;
  wire c105_d;
  wire c104_r;
  wire c104_a;
  wire c104_d;
  wire c103_r;
  wire c103_a;
  wire [16:0] c103_d;
  wire c102_r;
  wire c102_a;
  wire [16:0] c102_d;
  wire c101_r;
  wire c101_a;
  wire c100_r;
  wire c100_a;
  wire c99_r;
  wire c99_a;
  wire c98_r;
  wire c98_a;
  wire [16:0] c98_d;
  wire c97_r;
  wire c97_a;
  wire [16:0] c97_d;
  wire c96_r;
  wire c96_a;
  wire [15:0] c96_d;
  wire c95_r;
  wire c95_a;
  wire [17:0] c95_d;
  wire c94_r;
  wire c94_a;
  wire [16:0] c94_d;
  wire c93_r;
  wire c93_a;
  wire [16:0] c93_d;
  wire c92_r;
  wire c92_a;
  wire c92_d;
  wire c91_r;
  wire c91_a;
  wire [17:0] c91_d;
  wire c90_r;
  wire c90_a;
  wire [16:0] c90_d;
  wire c89_r;
  wire c89_a;
  wire [16:0] c89_d;
  wire c88_r;
  wire c88_a;
  wire c88_d;
  wire c87_r;
  wire c87_a;
  wire c87_d;
  wire c86_r;
  wire c86_a;
  wire c86_d;
  wire c85_r;
  wire c85_a;
  wire c85_d;
  wire c84_r;
  wire c84_a;
  wire [16:0] c84_d;
  wire c83_r;
  wire c83_a;
  wire [16:0] c83_d;
  wire c82_r;
  wire c82_a;
  wire c81_r;
  wire c81_a;
  wire c80_r;
  wire c80_a;
  wire c79_r;
  wire c79_a;
  wire [16:0] c79_d;
  wire c78_r;
  wire c78_a;
  wire [16:0] c78_d;
  wire c77_r;
  wire c77_a;
  wire [15:0] c77_d;
  wire c76_r;
  wire c76_a;
  wire [17:0] c76_d;
  wire c75_r;
  wire c75_a;
  wire [16:0] c75_d;
  wire c74_r;
  wire c74_a;
  wire [16:0] c74_d;
  wire c73_r;
  wire c73_a;
  wire c73_d;
  wire c72_r;
  wire c72_a;
  wire [17:0] c72_d;
  wire c71_r;
  wire c71_a;
  wire [16:0] c71_d;
  wire c70_r;
  wire c70_a;
  wire [16:0] c70_d;
  wire c69_r;
  wire c69_a;
  wire [16:0] c69_d;
  wire c68_r;
  wire c68_a;
  wire [16:0] c68_d;
  wire c67_r;
  wire c67_a;
  wire c66_r;
  wire c66_a;
  wire c65_r;
  wire c65_a;
  wire c64_r;
  wire c64_a;
  wire [16:0] c64_d;
  wire c63_r;
  wire c63_a;
  wire [16:0] c63_d;
  wire c62_r;
  wire c62_a;
  wire [15:0] c62_d;
  wire c61_r;
  wire c61_a;
  wire c61_d;
  wire c60_r;
  wire c60_a;
  wire c60_d;
  wire c59_r;
  wire c59_a;
  wire c59_d;
  wire c58_r;
  wire c58_a;
  wire c57_r;
  wire c57_a;
  wire c56_r;
  wire c56_a;
  wire c56_d;
  wire c55_r;
  wire c55_a;
  wire c54_r;
  wire c54_a;
  wire c54_d;
  wire c53_r;
  wire c53_a;
  wire c53_d;
  wire c52_r;
  wire c52_a;
  wire c52_d;
  wire c51_r;
  wire c51_a;
  wire c51_d;
  wire c50_r;
  wire c50_a;
  wire c50_d;
  wire c49_r;
  wire c49_a;
  wire [16:0] c49_d;
  wire c48_r;
  wire c48_a;
  wire [16:0] c48_d;
  wire c47_r;
  wire c47_a;
  wire c46_r;
  wire c46_a;
  wire c45_r;
  wire c45_a;
  wire c44_r;
  wire c44_a;
  wire [16:0] c44_d;
  wire c43_r;
  wire c43_a;
  wire [16:0] c43_d;
  wire c42_r;
  wire c42_a;
  wire [15:0] c42_d;
  wire c41_r;
  wire c41_a;
  wire [17:0] c41_d;
  wire c40_r;
  wire c40_a;
  wire [16:0] c40_d;
  wire c39_r;
  wire c39_a;
  wire [16:0] c39_d;
  wire c38_r;
  wire c38_a;
  wire c38_d;
  wire c37_r;
  wire c37_a;
  wire [17:0] c37_d;
  wire c36_r;
  wire c36_a;
  wire [16:0] c36_d;
  wire c35_r;
  wire c35_a;
  wire [16:0] c35_d;
  wire c34_r;
  wire c34_a;
  wire c34_d;
  wire c33_r;
  wire c33_a;
  wire c33_d;
  wire c32_r;
  wire c32_a;
  wire c32_d;
  wire c31_r;
  wire c31_a;
  wire c31_d;
  wire c30_r;
  wire c30_a;
  wire [16:0] c30_d;
  wire c29_r;
  wire c29_a;
  wire [16:0] c29_d;
  wire c28_r;
  wire c28_a;
  wire c27_r;
  wire c27_a;
  wire c26_r;
  wire c26_a;
  wire c25_r;
  wire c25_a;
  wire [16:0] c25_d;
  wire c24_r;
  wire c24_a;
  wire [16:0] c24_d;
  wire c23_r;
  wire c23_a;
  wire [15:0] c23_d;
  wire c22_r;
  wire c22_a;
  wire [17:0] c22_d;
  wire c21_r;
  wire c21_a;
  wire [16:0] c21_d;
  wire c20_r;
  wire c20_a;
  wire [16:0] c20_d;
  wire c19_r;
  wire c19_a;
  wire c19_d;
  wire c18_r;
  wire c18_a;
  wire [17:0] c18_d;
  wire c17_r;
  wire c17_a;
  wire [16:0] c17_d;
  wire c16_r;
  wire c16_a;
  wire [16:0] c16_d;
  wire c15_r;
  wire c15_a;
  wire [16:0] c15_d;
  wire c14_r;
  wire c14_a;
  wire [16:0] c14_d;
  wire c13_r;
  wire c13_a;
  wire c12_r;
  wire c12_a;
  wire c11_r;
  wire c11_a;
  wire c10_r;
  wire c10_a;
  wire [16:0] c10_d;
  wire c9_r;
  wire c9_a;
  wire [16:0] c9_d;
  wire c8_r;
  wire c8_a;
  wire [15:0] c8_d;
  wire c7_r;
  wire c7_a;
  wire c7_d;
  wire c6_r;
  wire c6_a;
  wire c5_r;
  wire c5_a;
  wire [15:0] c5_d;
  BrzVariable_8_2_s0_ I0 (c459_r, c459_a, c459_d, c451_r, c451_a, c451_d, c445_r, c445_a, c445_d);
  BrzVariable_8_1_s0_ I1 (c457_r, c457_a, c457_d, c439_r, c439_a, c439_d);
  BrzVariable_17_16_s0_ I2 (c454_r, c454_a, c454_d, c398_r, c398_a, c398_d, c394_r, c394_a, c394_d, c344_r, c344_a, c344_d, c340_r, c340_a, c340_d, c290_r, c290_a, c290_d, c286_r, c286_a, c286_d, c236_r, c236_a, c236_d, c232_r, c232_a, c232_d, c182_r, c182_a, c182_d, c178_r, c178_a, c178_d, c128_r, c128_a, c128_d, c124_r, c124_a, c124_d, c74_r, c74_a, c74_d, c70_r, c70_a, c70_d, c20_r, c20_a, c20_d, c16_r, c16_a,
		c16_d);
  BrzVariable_17_16_s0_ I3 (c449_r, c449_a, c449_d, c417_r, c417_a, c417_d, c413_r, c413_a, c413_d, c363_r, c363_a, c363_d, c359_r, c359_a, c359_d, c309_r, c309_a, c309_d, c305_r, c305_a, c305_d, c255_r, c255_a, c255_d, c251_r, c251_a, c251_d, c201_r, c201_a, c201_d, c197_r, c197_a, c197_d, c147_r, c147_a, c147_d, c143_r, c143_a, c143_d, c93_r, c93_a, c93_d, c89_r, c89_a, c89_d, c39_r, c39_a, c39_d, c35_r, c35_a,
		c35_d);
  BrzVariable_17_81_s657_1_2e_2e1_3b0_2e_2e0_m6m I4 (c463_r, c463_a, c463_d, c430_r, c430_a, c430_d, c428_r, c428_a, c428_d, c410_r, c410_a, c410_d, c409_r, c409_a, c409_d, c418_r, c418_a, c418_d, c414_r, c414_a, c414_d, c399_r, c399_a, c399_d, c395_r, c395_a, c395_d, c386_r, c386_a, c386_d, c385_r, c385_a, c385_d, c376_r, c376_a, c376_d, c374_r, c374_a, c374_d, c356_r, c356_a, c356_d, c355_r, c355_a, c355_d, c364_r, c364_a, c364_d, c360_r, c360_a,
		c360_d, c345_r, c345_a, c345_d, c341_r, c341_a, c341_d, c332_r, c332_a, c332_d, c331_r, c331_a, c331_d, c322_r, c322_a, c322_d, c320_r, c320_a, c320_d, c302_r, c302_a, c302_d, c301_r, c301_a, c301_d, c310_r, c310_a, c310_d, c306_r, c306_a, c306_d, c291_r, c291_a, c291_d, c287_r, c287_a, c287_d, c278_r, c278_a, c278_d, c277_r, c277_a, c277_d, c268_r, c268_a, c268_d, c266_r, c266_a, c266_d, c248_r, c248_a,
		c248_d, c247_r, c247_a, c247_d, c256_r, c256_a, c256_d, c252_r, c252_a, c252_d, c237_r, c237_a, c237_d, c233_r, c233_a, c233_d, c224_r, c224_a, c224_d, c223_r, c223_a, c223_d, c214_r, c214_a, c214_d, c212_r, c212_a, c212_d, c194_r, c194_a, c194_d, c193_r, c193_a, c193_d, c202_r, c202_a, c202_d, c198_r, c198_a, c198_d, c183_r, c183_a, c183_d, c179_r, c179_a, c179_d, c170_r, c170_a, c170_d, c169_r, c169_a,
		c169_d, c160_r, c160_a, c160_d, c158_r, c158_a, c158_d, c140_r, c140_a, c140_d, c139_r, c139_a, c139_d, c148_r, c148_a, c148_d, c144_r, c144_a, c144_d, c129_r, c129_a, c129_d, c125_r, c125_a, c125_d, c116_r, c116_a, c116_d, c115_r, c115_a, c115_d, c106_r, c106_a, c106_d, c104_r, c104_a, c104_d, c86_r, c86_a, c86_d, c85_r, c85_a, c85_d, c94_r, c94_a, c94_d, c90_r, c90_a, c90_d, c75_r, c75_a,
		c75_d, c71_r, c71_a, c71_d, c62_r, c62_a, c62_d, c61_r, c61_a, c61_d, c52_r, c52_a, c52_d, c50_r, c50_a, c50_d, c32_r, c32_a, c32_d, c31_r, c31_a, c31_d, c40_r, c40_a, c40_d, c36_r, c36_a, c36_d, c21_r, c21_a, c21_d, c17_r, c17_a, c17_d, c8_r, c8_a, c8_d, c7_r, c7_a, c7_d, c5_r, c5_a, c5_d);
  BrzCallMux_17_25 I5 (c10_r, c10_a, c10_d, c25_r, c25_a, c25_d, c44_r, c44_a, c44_d, c64_r, c64_a, c64_d, c79_r, c79_a, c79_d, c98_r, c98_a, c98_d, c118_r, c118_a, c118_d, c133_r, c133_a, c133_d, c152_r, c152_a, c152_d, c172_r, c172_a, c172_d, c187_r, c187_a, c187_d, c206_r, c206_a, c206_d, c226_r, c226_a, c226_d, c241_r, c241_a, c241_d, c260_r, c260_a, c260_d, c280_r, c280_a, c280_d, c295_r, c295_a,
		c295_d, c314_r, c314_a, c314_d, c334_r, c334_a, c334_d, c349_r, c349_a, c349_d, c368_r, c368_a, c368_d, c388_r, c388_a, c388_d, c403_r, c403_a, c403_d, c422_r, c422_a, c422_d, c443_r, c443_a, c443_d, c463_r, c463_a, c463_d);
  BrzLoop I6 (activate_0r, activate_0a, c462_r, c462_a);
  BrzSequence_19_s18_SSSSSSSSSSSSSSSSSS I7 (c462_r, c462_a, c461_r, c461_a, c456_r, c456_a, c435_r, c435_a, c436_r, c436_a, c381_r, c381_a, c382_r, c382_a, c327_r, c327_a, c328_r, c328_a, c273_r, c273_a, c274_r, c274_a, c219_r, c219_a, c220_r, c220_a, c165_r, c165_a, c166_r, c166_a, c111_r, c111_a, c112_r, c112_a, c57_r, c57_a, c58_r, c58_a, c6_r, c6_a);
  BrzConcur_2 I8 (c461_r, c461_a, c460_r, c460_a, c458_r, c458_a);
  BrzFetch_8_s5_false I9 (c460_r, c460_a, x_0r, x_0a, x_0d, c459_r, c459_a, c459_d);
  BrzFetch_8_s5_false I10 (c458_r, c458_a, y_0r, y_0a, y_0d, c457_r, c457_a, c457_d);
  BrzConcur_3 I11 (c456_r, c456_a, c455_r, c455_a, c450_r, c450_a, c444_r, c444_a);
  BrzFetch_17_s5_false I12 (c455_r, c455_a, c453_r, c453_a, c453_d, c454_r, c454_a, c454_d);
  BrzCombine_17_9_8 I13 (c453_r, c453_a, c453_d, c452_r, c452_a, c452_d, c451_r, c451_a, c451_d);
  BrzConstant_9_0 I14 (c452_r, c452_a, c452_d);
  BrzFetch_17_s5_false I15 (c450_r, c450_a, c448_r, c448_a, c448_d, c449_r, c449_a, c449_d);
  BrzCombine_17_9_8 I16 (c448_r, c448_a, c448_d, c447_r, c447_a, c447_d, c446_r, c446_a, c446_d);
  BrzConstant_9_0 I17 (c447_r, c447_a, c447_d);
  BrzUnaryFunc_8_8_s6_Negate_s4_true I18 (c446_r, c446_a, c446_d, c445_r, c445_a, c445_d);
  BrzFetch_17_s5_false I19 (c444_r, c444_a, c442_r, c442_a, c442_d, c443_r, c443_a, c443_d);
  BrzAdapt_17_9_s5_false_s5_false I20 (c442_r, c442_a, c442_d, c441_r, c441_a, c441_d);
  BrzCombine_9_1_8 I21 (c441_r, c441_a, c441_d, c440_r, c440_a, c440_d, c439_r, c439_a, c439_d);
  BrzConstant_1_0 I22 (c440_r, c440_a, c440_d);
  BrzCase_1_2_s5_0_3b1 I23 (c434_r, c434_a, c434_d, c389_r, c389_a, c433_r, c433_a);
  BrzFetch_1_s5_false I24 (c435_r, c435_a, c432_r, c432_a, c432_d, c437_r, c437_a, c437_d);
  BrzFetch_1_s5_false I25 (c436_r, c436_a, c438_r, c438_a, c438_d, c434_r, c434_a, c434_d);
  BrzVariable_1_1_s0_ I26 (c437_r, c437_a, c437_d, c438_r, c438_a, c438_d);
  BrzBar_2 I27 (c432_r, c432_a, c432_d, c433_r, c433_a, c412_r, c412_a, c412_d, c431_r, c431_a, c431_d, c404_r, c404_a, c423_r, c423_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I28 (c431_r, c431_a, c431_d, c430_r, c430_a, c430_d, c429_r, c429_a, c429_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I29 (c429_r, c429_a, c429_d, c428_r, c428_a, c428_d);
  BrzSequence_2_s1_S I30 (c423_r, c423_a, c424_r, c424_a, c425_r, c425_a);
  BrzFetch_17_s5_false I31 (c424_r, c424_a, c421_r, c421_a, c421_d, c426_r, c426_a, c426_d);
  BrzFetch_17_s5_false I32 (c425_r, c425_a, c427_r, c427_a, c427_d, c422_r, c422_a, c422_d);
  BrzVariable_17_1_s0_ I33 (c426_r, c426_a, c426_d, c427_r, c427_a, c427_d);
  BrzCombine_17_16_1 I34 (c421_r, c421_a, c421_d, c420_r, c420_a, c420_d, c416_r, c416_a, c416_d);
  BrzSlice_16_18_1 I35 (c420_r, c420_a, c420_d, c419_r, c419_a, c419_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I36 (c419_r, c419_a, c419_d, c418_r, c418_a, c418_d, c417_r, c417_a, c417_d);
  BrzSlice_1_18_16 I37 (c416_r, c416_a, c416_d, c415_r, c415_a, c415_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I38 (c415_r, c415_a, c415_d, c414_r, c414_a, c414_d, c413_r, c413_a, c413_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I39 (c412_r, c412_a, c412_d, c411_r, c411_a, c411_d, c409_r, c409_a, c409_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I40 (c411_r, c411_a, c411_d, c410_r, c410_a, c410_d);
  BrzSequence_2_s1_S I41 (c404_r, c404_a, c405_r, c405_a, c406_r, c406_a);
  BrzFetch_17_s5_false I42 (c405_r, c405_a, c402_r, c402_a, c402_d, c407_r, c407_a, c407_d);
  BrzFetch_17_s5_false I43 (c406_r, c406_a, c408_r, c408_a, c408_d, c403_r, c403_a, c403_d);
  BrzVariable_17_1_s0_ I44 (c407_r, c407_a, c407_d, c408_r, c408_a, c408_d);
  BrzCombine_17_16_1 I45 (c402_r, c402_a, c402_d, c401_r, c401_a, c401_d, c397_r, c397_a, c397_d);
  BrzSlice_16_18_1 I46 (c401_r, c401_a, c401_d, c400_r, c400_a, c400_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I47 (c400_r, c400_a, c400_d, c399_r, c399_a, c399_d, c398_r, c398_a, c398_d);
  BrzSlice_1_18_16 I48 (c397_r, c397_a, c397_d, c396_r, c396_a, c396_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I49 (c396_r, c396_a, c396_d, c395_r, c395_a, c395_d, c394_r, c394_a, c394_d);
  BrzSequence_2_s1_S I50 (c389_r, c389_a, c390_r, c390_a, c391_r, c391_a);
  BrzFetch_17_s5_false I51 (c390_r, c390_a, c387_r, c387_a, c387_d, c392_r, c392_a, c392_d);
  BrzFetch_17_s5_false I52 (c391_r, c391_a, c393_r, c393_a, c393_d, c388_r, c388_a, c388_d);
  BrzVariable_17_1_s0_ I53 (c392_r, c392_a, c392_d, c393_r, c393_a, c393_d);
  BrzCombine_17_16_1 I54 (c387_r, c387_a, c387_d, c386_r, c386_a, c386_d, c385_r, c385_a, c385_d);
  BrzCase_1_2_s5_0_3b1 I55 (c380_r, c380_a, c380_d, c335_r, c335_a, c379_r, c379_a);
  BrzFetch_1_s5_false I56 (c381_r, c381_a, c378_r, c378_a, c378_d, c383_r, c383_a, c383_d);
  BrzFetch_1_s5_false I57 (c382_r, c382_a, c384_r, c384_a, c384_d, c380_r, c380_a, c380_d);
  BrzVariable_1_1_s0_ I58 (c383_r, c383_a, c383_d, c384_r, c384_a, c384_d);
  BrzBar_2 I59 (c378_r, c378_a, c378_d, c379_r, c379_a, c358_r, c358_a, c358_d, c377_r, c377_a, c377_d, c350_r, c350_a, c369_r, c369_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I60 (c377_r, c377_a, c377_d, c376_r, c376_a, c376_d, c375_r, c375_a, c375_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I61 (c375_r, c375_a, c375_d, c374_r, c374_a, c374_d);
  BrzSequence_2_s1_S I62 (c369_r, c369_a, c370_r, c370_a, c371_r, c371_a);
  BrzFetch_17_s5_false I63 (c370_r, c370_a, c367_r, c367_a, c367_d, c372_r, c372_a, c372_d);
  BrzFetch_17_s5_false I64 (c371_r, c371_a, c373_r, c373_a, c373_d, c368_r, c368_a, c368_d);
  BrzVariable_17_1_s0_ I65 (c372_r, c372_a, c372_d, c373_r, c373_a, c373_d);
  BrzCombine_17_16_1 I66 (c367_r, c367_a, c367_d, c366_r, c366_a, c366_d, c362_r, c362_a, c362_d);
  BrzSlice_16_18_1 I67 (c366_r, c366_a, c366_d, c365_r, c365_a, c365_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I68 (c365_r, c365_a, c365_d, c364_r, c364_a, c364_d, c363_r, c363_a, c363_d);
  BrzSlice_1_18_16 I69 (c362_r, c362_a, c362_d, c361_r, c361_a, c361_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I70 (c361_r, c361_a, c361_d, c360_r, c360_a, c360_d, c359_r, c359_a, c359_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I71 (c358_r, c358_a, c358_d, c357_r, c357_a, c357_d, c355_r, c355_a, c355_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I72 (c357_r, c357_a, c357_d, c356_r, c356_a, c356_d);
  BrzSequence_2_s1_S I73 (c350_r, c350_a, c351_r, c351_a, c352_r, c352_a);
  BrzFetch_17_s5_false I74 (c351_r, c351_a, c348_r, c348_a, c348_d, c353_r, c353_a, c353_d);
  BrzFetch_17_s5_false I75 (c352_r, c352_a, c354_r, c354_a, c354_d, c349_r, c349_a, c349_d);
  BrzVariable_17_1_s0_ I76 (c353_r, c353_a, c353_d, c354_r, c354_a, c354_d);
  BrzCombine_17_16_1 I77 (c348_r, c348_a, c348_d, c347_r, c347_a, c347_d, c343_r, c343_a, c343_d);
  BrzSlice_16_18_1 I78 (c347_r, c347_a, c347_d, c346_r, c346_a, c346_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I79 (c346_r, c346_a, c346_d, c345_r, c345_a, c345_d, c344_r, c344_a, c344_d);
  BrzSlice_1_18_16 I80 (c343_r, c343_a, c343_d, c342_r, c342_a, c342_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I81 (c342_r, c342_a, c342_d, c341_r, c341_a, c341_d, c340_r, c340_a, c340_d);
  BrzSequence_2_s1_S I82 (c335_r, c335_a, c336_r, c336_a, c337_r, c337_a);
  BrzFetch_17_s5_false I83 (c336_r, c336_a, c333_r, c333_a, c333_d, c338_r, c338_a, c338_d);
  BrzFetch_17_s5_false I84 (c337_r, c337_a, c339_r, c339_a, c339_d, c334_r, c334_a, c334_d);
  BrzVariable_17_1_s0_ I85 (c338_r, c338_a, c338_d, c339_r, c339_a, c339_d);
  BrzCombine_17_16_1 I86 (c333_r, c333_a, c333_d, c332_r, c332_a, c332_d, c331_r, c331_a, c331_d);
  BrzCase_1_2_s5_0_3b1 I87 (c326_r, c326_a, c326_d, c281_r, c281_a, c325_r, c325_a);
  BrzFetch_1_s5_false I88 (c327_r, c327_a, c324_r, c324_a, c324_d, c329_r, c329_a, c329_d);
  BrzFetch_1_s5_false I89 (c328_r, c328_a, c330_r, c330_a, c330_d, c326_r, c326_a, c326_d);
  BrzVariable_1_1_s0_ I90 (c329_r, c329_a, c329_d, c330_r, c330_a, c330_d);
  BrzBar_2 I91 (c324_r, c324_a, c324_d, c325_r, c325_a, c304_r, c304_a, c304_d, c323_r, c323_a, c323_d, c296_r, c296_a, c315_r, c315_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I92 (c323_r, c323_a, c323_d, c322_r, c322_a, c322_d, c321_r, c321_a, c321_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I93 (c321_r, c321_a, c321_d, c320_r, c320_a, c320_d);
  BrzSequence_2_s1_S I94 (c315_r, c315_a, c316_r, c316_a, c317_r, c317_a);
  BrzFetch_17_s5_false I95 (c316_r, c316_a, c313_r, c313_a, c313_d, c318_r, c318_a, c318_d);
  BrzFetch_17_s5_false I96 (c317_r, c317_a, c319_r, c319_a, c319_d, c314_r, c314_a, c314_d);
  BrzVariable_17_1_s0_ I97 (c318_r, c318_a, c318_d, c319_r, c319_a, c319_d);
  BrzCombine_17_16_1 I98 (c313_r, c313_a, c313_d, c312_r, c312_a, c312_d, c308_r, c308_a, c308_d);
  BrzSlice_16_18_1 I99 (c312_r, c312_a, c312_d, c311_r, c311_a, c311_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I100 (c311_r, c311_a, c311_d, c310_r, c310_a, c310_d, c309_r, c309_a, c309_d);
  BrzSlice_1_18_16 I101 (c308_r, c308_a, c308_d, c307_r, c307_a, c307_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I102 (c307_r, c307_a, c307_d, c306_r, c306_a, c306_d, c305_r, c305_a, c305_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I103 (c304_r, c304_a, c304_d, c303_r, c303_a, c303_d, c301_r, c301_a, c301_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I104 (c303_r, c303_a, c303_d, c302_r, c302_a, c302_d);
  BrzSequence_2_s1_S I105 (c296_r, c296_a, c297_r, c297_a, c298_r, c298_a);
  BrzFetch_17_s5_false I106 (c297_r, c297_a, c294_r, c294_a, c294_d, c299_r, c299_a, c299_d);
  BrzFetch_17_s5_false I107 (c298_r, c298_a, c300_r, c300_a, c300_d, c295_r, c295_a, c295_d);
  BrzVariable_17_1_s0_ I108 (c299_r, c299_a, c299_d, c300_r, c300_a, c300_d);
  BrzCombine_17_16_1 I109 (c294_r, c294_a, c294_d, c293_r, c293_a, c293_d, c289_r, c289_a, c289_d);
  BrzSlice_16_18_1 I110 (c293_r, c293_a, c293_d, c292_r, c292_a, c292_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I111 (c292_r, c292_a, c292_d, c291_r, c291_a, c291_d, c290_r, c290_a, c290_d);
  BrzSlice_1_18_16 I112 (c289_r, c289_a, c289_d, c288_r, c288_a, c288_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I113 (c288_r, c288_a, c288_d, c287_r, c287_a, c287_d, c286_r, c286_a, c286_d);
  BrzSequence_2_s1_S I114 (c281_r, c281_a, c282_r, c282_a, c283_r, c283_a);
  BrzFetch_17_s5_false I115 (c282_r, c282_a, c279_r, c279_a, c279_d, c284_r, c284_a, c284_d);
  BrzFetch_17_s5_false I116 (c283_r, c283_a, c285_r, c285_a, c285_d, c280_r, c280_a, c280_d);
  BrzVariable_17_1_s0_ I117 (c284_r, c284_a, c284_d, c285_r, c285_a, c285_d);
  BrzCombine_17_16_1 I118 (c279_r, c279_a, c279_d, c278_r, c278_a, c278_d, c277_r, c277_a, c277_d);
  BrzCase_1_2_s5_0_3b1 I119 (c272_r, c272_a, c272_d, c227_r, c227_a, c271_r, c271_a);
  BrzFetch_1_s5_false I120 (c273_r, c273_a, c270_r, c270_a, c270_d, c275_r, c275_a, c275_d);
  BrzFetch_1_s5_false I121 (c274_r, c274_a, c276_r, c276_a, c276_d, c272_r, c272_a, c272_d);
  BrzVariable_1_1_s0_ I122 (c275_r, c275_a, c275_d, c276_r, c276_a, c276_d);
  BrzBar_2 I123 (c270_r, c270_a, c270_d, c271_r, c271_a, c250_r, c250_a, c250_d, c269_r, c269_a, c269_d, c242_r, c242_a, c261_r, c261_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I124 (c269_r, c269_a, c269_d, c268_r, c268_a, c268_d, c267_r, c267_a, c267_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I125 (c267_r, c267_a, c267_d, c266_r, c266_a, c266_d);
  BrzSequence_2_s1_S I126 (c261_r, c261_a, c262_r, c262_a, c263_r, c263_a);
  BrzFetch_17_s5_false I127 (c262_r, c262_a, c259_r, c259_a, c259_d, c264_r, c264_a, c264_d);
  BrzFetch_17_s5_false I128 (c263_r, c263_a, c265_r, c265_a, c265_d, c260_r, c260_a, c260_d);
  BrzVariable_17_1_s0_ I129 (c264_r, c264_a, c264_d, c265_r, c265_a, c265_d);
  BrzCombine_17_16_1 I130 (c259_r, c259_a, c259_d, c258_r, c258_a, c258_d, c254_r, c254_a, c254_d);
  BrzSlice_16_18_1 I131 (c258_r, c258_a, c258_d, c257_r, c257_a, c257_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I132 (c257_r, c257_a, c257_d, c256_r, c256_a, c256_d, c255_r, c255_a, c255_d);
  BrzSlice_1_18_16 I133 (c254_r, c254_a, c254_d, c253_r, c253_a, c253_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I134 (c253_r, c253_a, c253_d, c252_r, c252_a, c252_d, c251_r, c251_a, c251_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I135 (c250_r, c250_a, c250_d, c249_r, c249_a, c249_d, c247_r, c247_a, c247_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I136 (c249_r, c249_a, c249_d, c248_r, c248_a, c248_d);
  BrzSequence_2_s1_S I137 (c242_r, c242_a, c243_r, c243_a, c244_r, c244_a);
  BrzFetch_17_s5_false I138 (c243_r, c243_a, c240_r, c240_a, c240_d, c245_r, c245_a, c245_d);
  BrzFetch_17_s5_false I139 (c244_r, c244_a, c246_r, c246_a, c246_d, c241_r, c241_a, c241_d);
  BrzVariable_17_1_s0_ I140 (c245_r, c245_a, c245_d, c246_r, c246_a, c246_d);
  BrzCombine_17_16_1 I141 (c240_r, c240_a, c240_d, c239_r, c239_a, c239_d, c235_r, c235_a, c235_d);
  BrzSlice_16_18_1 I142 (c239_r, c239_a, c239_d, c238_r, c238_a, c238_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I143 (c238_r, c238_a, c238_d, c237_r, c237_a, c237_d, c236_r, c236_a, c236_d);
  BrzSlice_1_18_16 I144 (c235_r, c235_a, c235_d, c234_r, c234_a, c234_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I145 (c234_r, c234_a, c234_d, c233_r, c233_a, c233_d, c232_r, c232_a, c232_d);
  BrzSequence_2_s1_S I146 (c227_r, c227_a, c228_r, c228_a, c229_r, c229_a);
  BrzFetch_17_s5_false I147 (c228_r, c228_a, c225_r, c225_a, c225_d, c230_r, c230_a, c230_d);
  BrzFetch_17_s5_false I148 (c229_r, c229_a, c231_r, c231_a, c231_d, c226_r, c226_a, c226_d);
  BrzVariable_17_1_s0_ I149 (c230_r, c230_a, c230_d, c231_r, c231_a, c231_d);
  BrzCombine_17_16_1 I150 (c225_r, c225_a, c225_d, c224_r, c224_a, c224_d, c223_r, c223_a, c223_d);
  BrzCase_1_2_s5_0_3b1 I151 (c218_r, c218_a, c218_d, c173_r, c173_a, c217_r, c217_a);
  BrzFetch_1_s5_false I152 (c219_r, c219_a, c216_r, c216_a, c216_d, c221_r, c221_a, c221_d);
  BrzFetch_1_s5_false I153 (c220_r, c220_a, c222_r, c222_a, c222_d, c218_r, c218_a, c218_d);
  BrzVariable_1_1_s0_ I154 (c221_r, c221_a, c221_d, c222_r, c222_a, c222_d);
  BrzBar_2 I155 (c216_r, c216_a, c216_d, c217_r, c217_a, c196_r, c196_a, c196_d, c215_r, c215_a, c215_d, c188_r, c188_a, c207_r, c207_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I156 (c215_r, c215_a, c215_d, c214_r, c214_a, c214_d, c213_r, c213_a, c213_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I157 (c213_r, c213_a, c213_d, c212_r, c212_a, c212_d);
  BrzSequence_2_s1_S I158 (c207_r, c207_a, c208_r, c208_a, c209_r, c209_a);
  BrzFetch_17_s5_false I159 (c208_r, c208_a, c205_r, c205_a, c205_d, c210_r, c210_a, c210_d);
  BrzFetch_17_s5_false I160 (c209_r, c209_a, c211_r, c211_a, c211_d, c206_r, c206_a, c206_d);
  BrzVariable_17_1_s0_ I161 (c210_r, c210_a, c210_d, c211_r, c211_a, c211_d);
  BrzCombine_17_16_1 I162 (c205_r, c205_a, c205_d, c204_r, c204_a, c204_d, c200_r, c200_a, c200_d);
  BrzSlice_16_18_1 I163 (c204_r, c204_a, c204_d, c203_r, c203_a, c203_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I164 (c203_r, c203_a, c203_d, c202_r, c202_a, c202_d, c201_r, c201_a, c201_d);
  BrzSlice_1_18_16 I165 (c200_r, c200_a, c200_d, c199_r, c199_a, c199_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I166 (c199_r, c199_a, c199_d, c198_r, c198_a, c198_d, c197_r, c197_a, c197_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I167 (c196_r, c196_a, c196_d, c195_r, c195_a, c195_d, c193_r, c193_a, c193_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I168 (c195_r, c195_a, c195_d, c194_r, c194_a, c194_d);
  BrzSequence_2_s1_S I169 (c188_r, c188_a, c189_r, c189_a, c190_r, c190_a);
  BrzFetch_17_s5_false I170 (c189_r, c189_a, c186_r, c186_a, c186_d, c191_r, c191_a, c191_d);
  BrzFetch_17_s5_false I171 (c190_r, c190_a, c192_r, c192_a, c192_d, c187_r, c187_a, c187_d);
  BrzVariable_17_1_s0_ I172 (c191_r, c191_a, c191_d, c192_r, c192_a, c192_d);
  BrzCombine_17_16_1 I173 (c186_r, c186_a, c186_d, c185_r, c185_a, c185_d, c181_r, c181_a, c181_d);
  BrzSlice_16_18_1 I174 (c185_r, c185_a, c185_d, c184_r, c184_a, c184_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I175 (c184_r, c184_a, c184_d, c183_r, c183_a, c183_d, c182_r, c182_a, c182_d);
  BrzSlice_1_18_16 I176 (c181_r, c181_a, c181_d, c180_r, c180_a, c180_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I177 (c180_r, c180_a, c180_d, c179_r, c179_a, c179_d, c178_r, c178_a, c178_d);
  BrzSequence_2_s1_S I178 (c173_r, c173_a, c174_r, c174_a, c175_r, c175_a);
  BrzFetch_17_s5_false I179 (c174_r, c174_a, c171_r, c171_a, c171_d, c176_r, c176_a, c176_d);
  BrzFetch_17_s5_false I180 (c175_r, c175_a, c177_r, c177_a, c177_d, c172_r, c172_a, c172_d);
  BrzVariable_17_1_s0_ I181 (c176_r, c176_a, c176_d, c177_r, c177_a, c177_d);
  BrzCombine_17_16_1 I182 (c171_r, c171_a, c171_d, c170_r, c170_a, c170_d, c169_r, c169_a, c169_d);
  BrzCase_1_2_s5_0_3b1 I183 (c164_r, c164_a, c164_d, c119_r, c119_a, c163_r, c163_a);
  BrzFetch_1_s5_false I184 (c165_r, c165_a, c162_r, c162_a, c162_d, c167_r, c167_a, c167_d);
  BrzFetch_1_s5_false I185 (c166_r, c166_a, c168_r, c168_a, c168_d, c164_r, c164_a, c164_d);
  BrzVariable_1_1_s0_ I186 (c167_r, c167_a, c167_d, c168_r, c168_a, c168_d);
  BrzBar_2 I187 (c162_r, c162_a, c162_d, c163_r, c163_a, c142_r, c142_a, c142_d, c161_r, c161_a, c161_d, c134_r, c134_a, c153_r, c153_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I188 (c161_r, c161_a, c161_d, c160_r, c160_a, c160_d, c159_r, c159_a, c159_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I189 (c159_r, c159_a, c159_d, c158_r, c158_a, c158_d);
  BrzSequence_2_s1_S I190 (c153_r, c153_a, c154_r, c154_a, c155_r, c155_a);
  BrzFetch_17_s5_false I191 (c154_r, c154_a, c151_r, c151_a, c151_d, c156_r, c156_a, c156_d);
  BrzFetch_17_s5_false I192 (c155_r, c155_a, c157_r, c157_a, c157_d, c152_r, c152_a, c152_d);
  BrzVariable_17_1_s0_ I193 (c156_r, c156_a, c156_d, c157_r, c157_a, c157_d);
  BrzCombine_17_16_1 I194 (c151_r, c151_a, c151_d, c150_r, c150_a, c150_d, c146_r, c146_a, c146_d);
  BrzSlice_16_18_1 I195 (c150_r, c150_a, c150_d, c149_r, c149_a, c149_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I196 (c149_r, c149_a, c149_d, c148_r, c148_a, c148_d, c147_r, c147_a, c147_d);
  BrzSlice_1_18_16 I197 (c146_r, c146_a, c146_d, c145_r, c145_a, c145_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I198 (c145_r, c145_a, c145_d, c144_r, c144_a, c144_d, c143_r, c143_a, c143_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I199 (c142_r, c142_a, c142_d, c141_r, c141_a, c141_d, c139_r, c139_a, c139_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I200 (c141_r, c141_a, c141_d, c140_r, c140_a, c140_d);
  BrzSequence_2_s1_S I201 (c134_r, c134_a, c135_r, c135_a, c136_r, c136_a);
  BrzFetch_17_s5_false I202 (c135_r, c135_a, c132_r, c132_a, c132_d, c137_r, c137_a, c137_d);
  BrzFetch_17_s5_false I203 (c136_r, c136_a, c138_r, c138_a, c138_d, c133_r, c133_a, c133_d);
  BrzVariable_17_1_s0_ I204 (c137_r, c137_a, c137_d, c138_r, c138_a, c138_d);
  BrzCombine_17_16_1 I205 (c132_r, c132_a, c132_d, c131_r, c131_a, c131_d, c127_r, c127_a, c127_d);
  BrzSlice_16_18_1 I206 (c131_r, c131_a, c131_d, c130_r, c130_a, c130_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I207 (c130_r, c130_a, c130_d, c129_r, c129_a, c129_d, c128_r, c128_a, c128_d);
  BrzSlice_1_18_16 I208 (c127_r, c127_a, c127_d, c126_r, c126_a, c126_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I209 (c126_r, c126_a, c126_d, c125_r, c125_a, c125_d, c124_r, c124_a, c124_d);
  BrzSequence_2_s1_S I210 (c119_r, c119_a, c120_r, c120_a, c121_r, c121_a);
  BrzFetch_17_s5_false I211 (c120_r, c120_a, c117_r, c117_a, c117_d, c122_r, c122_a, c122_d);
  BrzFetch_17_s5_false I212 (c121_r, c121_a, c123_r, c123_a, c123_d, c118_r, c118_a, c118_d);
  BrzVariable_17_1_s0_ I213 (c122_r, c122_a, c122_d, c123_r, c123_a, c123_d);
  BrzCombine_17_16_1 I214 (c117_r, c117_a, c117_d, c116_r, c116_a, c116_d, c115_r, c115_a, c115_d);
  BrzCase_1_2_s5_0_3b1 I215 (c110_r, c110_a, c110_d, c65_r, c65_a, c109_r, c109_a);
  BrzFetch_1_s5_false I216 (c111_r, c111_a, c108_r, c108_a, c108_d, c113_r, c113_a, c113_d);
  BrzFetch_1_s5_false I217 (c112_r, c112_a, c114_r, c114_a, c114_d, c110_r, c110_a, c110_d);
  BrzVariable_1_1_s0_ I218 (c113_r, c113_a, c113_d, c114_r, c114_a, c114_d);
  BrzBar_2 I219 (c108_r, c108_a, c108_d, c109_r, c109_a, c88_r, c88_a, c88_d, c107_r, c107_a, c107_d, c80_r, c80_a, c99_r, c99_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I220 (c107_r, c107_a, c107_d, c106_r, c106_a, c106_d, c105_r, c105_a, c105_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I221 (c105_r, c105_a, c105_d, c104_r, c104_a, c104_d);
  BrzSequence_2_s1_S I222 (c99_r, c99_a, c100_r, c100_a, c101_r, c101_a);
  BrzFetch_17_s5_false I223 (c100_r, c100_a, c97_r, c97_a, c97_d, c102_r, c102_a, c102_d);
  BrzFetch_17_s5_false I224 (c101_r, c101_a, c103_r, c103_a, c103_d, c98_r, c98_a, c98_d);
  BrzVariable_17_1_s0_ I225 (c102_r, c102_a, c102_d, c103_r, c103_a, c103_d);
  BrzCombine_17_16_1 I226 (c97_r, c97_a, c97_d, c96_r, c96_a, c96_d, c92_r, c92_a, c92_d);
  BrzSlice_16_18_1 I227 (c96_r, c96_a, c96_d, c95_r, c95_a, c95_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I228 (c95_r, c95_a, c95_d, c94_r, c94_a, c94_d, c93_r, c93_a, c93_d);
  BrzSlice_1_18_16 I229 (c92_r, c92_a, c92_d, c91_r, c91_a, c91_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I230 (c91_r, c91_a, c91_d, c90_r, c90_a, c90_d, c89_r, c89_a, c89_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I231 (c88_r, c88_a, c88_d, c87_r, c87_a, c87_d, c85_r, c85_a, c85_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I232 (c87_r, c87_a, c87_d, c86_r, c86_a, c86_d);
  BrzSequence_2_s1_S I233 (c80_r, c80_a, c81_r, c81_a, c82_r, c82_a);
  BrzFetch_17_s5_false I234 (c81_r, c81_a, c78_r, c78_a, c78_d, c83_r, c83_a, c83_d);
  BrzFetch_17_s5_false I235 (c82_r, c82_a, c84_r, c84_a, c84_d, c79_r, c79_a, c79_d);
  BrzVariable_17_1_s0_ I236 (c83_r, c83_a, c83_d, c84_r, c84_a, c84_d);
  BrzCombine_17_16_1 I237 (c78_r, c78_a, c78_d, c77_r, c77_a, c77_d, c73_r, c73_a, c73_d);
  BrzSlice_16_18_1 I238 (c77_r, c77_a, c77_d, c76_r, c76_a, c76_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I239 (c76_r, c76_a, c76_d, c75_r, c75_a, c75_d, c74_r, c74_a, c74_d);
  BrzSlice_1_18_16 I240 (c73_r, c73_a, c73_d, c72_r, c72_a, c72_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I241 (c72_r, c72_a, c72_d, c71_r, c71_a, c71_d, c70_r, c70_a, c70_d);
  BrzSequence_2_s1_S I242 (c65_r, c65_a, c66_r, c66_a, c67_r, c67_a);
  BrzFetch_17_s5_false I243 (c66_r, c66_a, c63_r, c63_a, c63_d, c68_r, c68_a, c68_d);
  BrzFetch_17_s5_false I244 (c67_r, c67_a, c69_r, c69_a, c69_d, c64_r, c64_a, c64_d);
  BrzVariable_17_1_s0_ I245 (c68_r, c68_a, c68_d, c69_r, c69_a, c69_d);
  BrzCombine_17_16_1 I246 (c63_r, c63_a, c63_d, c62_r, c62_a, c62_d, c61_r, c61_a, c61_d);
  BrzCase_1_2_s5_0_3b1 I247 (c56_r, c56_a, c56_d, c11_r, c11_a, c55_r, c55_a);
  BrzFetch_1_s5_false I248 (c57_r, c57_a, c54_r, c54_a, c54_d, c59_r, c59_a, c59_d);
  BrzFetch_1_s5_false I249 (c58_r, c58_a, c60_r, c60_a, c60_d, c56_r, c56_a, c56_d);
  BrzVariable_1_1_s0_ I250 (c59_r, c59_a, c59_d, c60_r, c60_a, c60_d);
  BrzBar_2 I251 (c54_r, c54_a, c54_d, c55_r, c55_a, c34_r, c34_a, c34_d, c53_r, c53_a, c53_d, c26_r, c26_a, c45_r, c45_a);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I252 (c53_r, c53_a, c53_d, c52_r, c52_a, c52_d, c51_r, c51_a, c51_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I253 (c51_r, c51_a, c51_d, c50_r, c50_a, c50_d);
  BrzSequence_2_s1_S I254 (c45_r, c45_a, c46_r, c46_a, c47_r, c47_a);
  BrzFetch_17_s5_false I255 (c46_r, c46_a, c43_r, c43_a, c43_d, c48_r, c48_a, c48_d);
  BrzFetch_17_s5_false I256 (c47_r, c47_a, c49_r, c49_a, c49_d, c44_r, c44_a, c44_d);
  BrzVariable_17_1_s0_ I257 (c48_r, c48_a, c48_d, c49_r, c49_a, c49_d);
  BrzCombine_17_16_1 I258 (c43_r, c43_a, c43_d, c42_r, c42_a, c42_d, c38_r, c38_a, c38_d);
  BrzSlice_16_18_1 I259 (c42_r, c42_a, c42_d, c41_r, c41_a, c41_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I260 (c41_r, c41_a, c41_d, c40_r, c40_a, c40_d, c39_r, c39_a, c39_d);
  BrzSlice_1_18_16 I261 (c38_r, c38_a, c38_d, c37_r, c37_a, c37_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I262 (c37_r, c37_a, c37_d, c36_r, c36_a, c36_d, c35_r, c35_a, c35_d);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m1m I263 (c34_r, c34_a, c34_d, c33_r, c33_a, c33_d, c31_r, c31_a, c31_d);
  BrzUnaryFunc_1_1_s6_Invert_s5_false I264 (c33_r, c33_a, c33_d, c32_r, c32_a, c32_d);
  BrzSequence_2_s1_S I265 (c26_r, c26_a, c27_r, c27_a, c28_r, c28_a);
  BrzFetch_17_s5_false I266 (c27_r, c27_a, c24_r, c24_a, c24_d, c29_r, c29_a, c29_d);
  BrzFetch_17_s5_false I267 (c28_r, c28_a, c30_r, c30_a, c30_d, c25_r, c25_a, c25_d);
  BrzVariable_17_1_s0_ I268 (c29_r, c29_a, c29_d, c30_r, c30_a, c30_d);
  BrzCombine_17_16_1 I269 (c24_r, c24_a, c24_d, c23_r, c23_a, c23_d, c19_r, c19_a, c19_d);
  BrzSlice_16_18_1 I270 (c23_r, c23_a, c23_d, c22_r, c22_a, c22_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I271 (c22_r, c22_a, c22_d, c21_r, c21_a, c21_d, c20_r, c20_a, c20_d);
  BrzSlice_1_18_16 I272 (c19_r, c19_a, c19_d, c18_r, c18_a, c18_d);
  BrzBinaryFunc_18_17_17_s3_Add_s4_true_s4_t_m5m I273 (c18_r, c18_a, c18_d, c17_r, c17_a, c17_d, c16_r, c16_a, c16_d);
  BrzSequence_2_s1_S I274 (c11_r, c11_a, c12_r, c12_a, c13_r, c13_a);
  BrzFetch_17_s5_false I275 (c12_r, c12_a, c9_r, c9_a, c9_d, c14_r, c14_a, c14_d);
  BrzFetch_17_s5_false I276 (c13_r, c13_a, c15_r, c15_a, c15_d, c10_r, c10_a, c10_d);
  BrzVariable_17_1_s0_ I277 (c14_r, c14_a, c14_d, c15_r, c15_a, c15_d);
  BrzCombine_17_16_1 I278 (c9_r, c9_a, c9_d, c8_r, c8_a, c8_d, c7_r, c7_a, c7_d);
  BrzFetch_16_s5_false I279 (c6_r, c6_a, c5_r, c5_a, c5_d, z_0r, z_0a, z_0d);
endmodule

